module cpu (clk, reset, DI, IRQ, NMI, RDY, AB, DO, WE);

input clk;
input reset;
input IRQ;
input NMI;
input RDY;
output WE;
input [7:0] DI;
output [15:0] AB;
output [7:0] DO;

wire vdd = 1'b1;
wire gnd = 1'b0;

	BUFX4 BUFX4_1 ( .A(_1466_), .Y(_1466__bF_buf4) );
	BUFX4 BUFX4_2 ( .A(_1466_), .Y(_1466__bF_buf3) );
	BUFX4 BUFX4_3 ( .A(_1466_), .Y(_1466__bF_buf2) );
	BUFX4 BUFX4_4 ( .A(_1466_), .Y(_1466__bF_buf1) );
	BUFX4 BUFX4_5 ( .A(_1466_), .Y(_1466__bF_buf0) );
	BUFX4 BUFX4_6 ( .A(clk), .Y(clk_bF_buf11) );
	BUFX4 BUFX4_7 ( .A(clk), .Y(clk_bF_buf10) );
	BUFX4 BUFX4_8 ( .A(clk), .Y(clk_bF_buf9) );
	BUFX4 BUFX4_9 ( .A(clk), .Y(clk_bF_buf8) );
	BUFX4 BUFX4_10 ( .A(clk), .Y(clk_bF_buf7) );
	BUFX4 BUFX4_11 ( .A(clk), .Y(clk_bF_buf6) );
	BUFX4 BUFX4_12 ( .A(clk), .Y(clk_bF_buf5) );
	BUFX4 BUFX4_13 ( .A(clk), .Y(clk_bF_buf4) );
	BUFX4 BUFX4_14 ( .A(clk), .Y(clk_bF_buf3) );
	BUFX4 BUFX4_15 ( .A(clk), .Y(clk_bF_buf2) );
	BUFX4 BUFX4_16 ( .A(clk), .Y(clk_bF_buf1) );
	BUFX4 BUFX4_17 ( .A(clk), .Y(clk_bF_buf0) );
	BUFX4 BUFX4_18 ( .A(_936_), .Y(_936__bF_buf3) );
	BUFX4 BUFX4_19 ( .A(_936_), .Y(_936__bF_buf2) );
	BUFX2 BUFX2_1 ( .A(_936_), .Y(_936__bF_buf1) );
	BUFX4 BUFX4_20 ( .A(_936_), .Y(_936__bF_buf0) );
	BUFX4 BUFX4_21 ( .A(_882_), .Y(_882__bF_buf5) );
	BUFX4 BUFX4_22 ( .A(_882_), .Y(_882__bF_buf4) );
	BUFX4 BUFX4_23 ( .A(_882_), .Y(_882__bF_buf3) );
	BUFX4 BUFX4_24 ( .A(_882_), .Y(_882__bF_buf2) );
	BUFX4 BUFX4_25 ( .A(_882_), .Y(_882__bF_buf1) );
	BUFX4 BUFX4_26 ( .A(_882_), .Y(_882__bF_buf0) );
	BUFX2 BUFX2_2 ( .A(_1717_), .Y(_1717__bF_buf3) );
	BUFX4 BUFX4_27 ( .A(_1717_), .Y(_1717__bF_buf2) );
	BUFX4 BUFX4_28 ( .A(_1717_), .Y(_1717__bF_buf1) );
	BUFX4 BUFX4_29 ( .A(_1717_), .Y(_1717__bF_buf0) );
	BUFX4 BUFX4_30 ( .A(_886_), .Y(_886__bF_buf4) );
	BUFX4 BUFX4_31 ( .A(_886_), .Y(_886__bF_buf3) );
	BUFX4 BUFX4_32 ( .A(_886_), .Y(_886__bF_buf2) );
	BUFX4 BUFX4_33 ( .A(_886_), .Y(_886__bF_buf1) );
	BUFX4 BUFX4_34 ( .A(_886_), .Y(_886__bF_buf0) );
	BUFX4 BUFX4_35 ( .A(_881_), .Y(_881__bF_buf7) );
	BUFX4 BUFX4_36 ( .A(_881_), .Y(_881__bF_buf6) );
	BUFX4 BUFX4_37 ( .A(_881_), .Y(_881__bF_buf5) );
	BUFX4 BUFX4_38 ( .A(_881_), .Y(_881__bF_buf4) );
	BUFX4 BUFX4_39 ( .A(_881_), .Y(_881__bF_buf3) );
	BUFX4 BUFX4_40 ( .A(_881_), .Y(_881__bF_buf2) );
	BUFX4 BUFX4_41 ( .A(_881_), .Y(_881__bF_buf1) );
	BUFX4 BUFX4_42 ( .A(_881_), .Y(_881__bF_buf0) );
	BUFX4 BUFX4_43 ( .A(RDY), .Y(RDY_bF_buf8) );
	BUFX4 BUFX4_44 ( .A(RDY), .Y(RDY_bF_buf7) );
	BUFX4 BUFX4_45 ( .A(RDY), .Y(RDY_bF_buf6) );
	BUFX4 BUFX4_46 ( .A(RDY), .Y(RDY_bF_buf5) );
	BUFX4 BUFX4_47 ( .A(RDY), .Y(RDY_bF_buf4) );
	BUFX4 BUFX4_48 ( .A(RDY), .Y(RDY_bF_buf3) );
	BUFX4 BUFX4_49 ( .A(RDY), .Y(RDY_bF_buf2) );
	BUFX4 BUFX4_50 ( .A(RDY), .Y(RDY_bF_buf1) );
	BUFX4 BUFX4_51 ( .A(RDY), .Y(RDY_bF_buf0) );
	BUFX4 BUFX4_52 ( .A(_957_), .Y(_957__bF_buf4) );
	BUFX4 BUFX4_53 ( .A(_957_), .Y(_957__bF_buf3) );
	BUFX4 BUFX4_54 ( .A(_957_), .Y(_957__bF_buf2) );
	BUFX4 BUFX4_55 ( .A(_957_), .Y(_957__bF_buf1) );
	BUFX4 BUFX4_56 ( .A(_957_), .Y(_957__bF_buf0) );
	BUFX4 BUFX4_57 ( .A(_885_), .Y(_885__bF_buf4) );
	BUFX4 BUFX4_58 ( .A(_885_), .Y(_885__bF_buf3) );
	BUFX4 BUFX4_59 ( .A(_885_), .Y(_885__bF_buf2) );
	BUFX4 BUFX4_60 ( .A(_885_), .Y(_885__bF_buf1) );
	BUFX4 BUFX4_61 ( .A(_885_), .Y(_885__bF_buf0) );
	BUFX4 BUFX4_62 ( .A(_910_), .Y(_910__bF_buf4) );
	BUFX4 BUFX4_63 ( .A(_910_), .Y(_910__bF_buf3) );
	BUFX4 BUFX4_64 ( .A(_910_), .Y(_910__bF_buf2) );
	BUFX4 BUFX4_65 ( .A(_910_), .Y(_910__bF_buf1) );
	BUFX4 BUFX4_66 ( .A(_910_), .Y(_910__bF_buf0) );
	BUFX2 BUFX2_3 ( .A(_896_), .Y(_896__bF_buf3) );
	BUFX2 BUFX2_4 ( .A(_896_), .Y(_896__bF_buf2) );
	BUFX2 BUFX2_5 ( .A(_896_), .Y(_896__bF_buf1) );
	BUFX2 BUFX2_6 ( .A(_896_), .Y(_896__bF_buf0) );
	BUFX4 BUFX4_67 ( .A(_535_), .Y(_535__bF_buf4) );
	BUFX4 BUFX4_68 ( .A(_535_), .Y(_535__bF_buf3) );
	BUFX4 BUFX4_69 ( .A(_535_), .Y(_535__bF_buf2) );
	BUFX4 BUFX4_70 ( .A(_535_), .Y(_535__bF_buf1) );
	BUFX4 BUFX4_71 ( .A(_535_), .Y(_535__bF_buf0) );
	BUFX4 BUFX4_72 ( .A(_1034_), .Y(_1034__bF_buf3) );
	BUFX4 BUFX4_73 ( .A(_1034_), .Y(_1034__bF_buf2) );
	BUFX2 BUFX2_7 ( .A(_1034_), .Y(_1034__bF_buf1) );
	BUFX2 BUFX2_8 ( .A(_1034_), .Y(_1034__bF_buf0) );
	BUFX4 BUFX4_74 ( .A(_1057_), .Y(_1057__bF_buf3) );
	BUFX4 BUFX4_75 ( .A(_1057_), .Y(_1057__bF_buf2) );
	BUFX4 BUFX4_76 ( .A(_1057_), .Y(_1057__bF_buf1) );
	BUFX4 BUFX4_77 ( .A(_1057_), .Y(_1057__bF_buf0) );
	BUFX4 BUFX4_78 ( .A(_1022_), .Y(_1022__bF_buf3) );
	BUFX4 BUFX4_79 ( .A(_1022_), .Y(_1022__bF_buf2) );
	BUFX4 BUFX4_80 ( .A(_1022_), .Y(_1022__bF_buf1) );
	BUFX4 BUFX4_81 ( .A(_1022_), .Y(_1022__bF_buf0) );
	BUFX4 BUFX4_82 ( .A(_937_), .Y(_937__bF_buf4) );
	BUFX4 BUFX4_83 ( .A(_937_), .Y(_937__bF_buf3) );
	BUFX4 BUFX4_84 ( .A(_937_), .Y(_937__bF_buf2) );
	BUFX4 BUFX4_85 ( .A(_937_), .Y(_937__bF_buf1) );
	BUFX4 BUFX4_86 ( .A(_937_), .Y(_937__bF_buf0) );
	BUFX4 BUFX4_87 ( .A(_962_), .Y(_962__bF_buf4) );
	BUFX4 BUFX4_88 ( .A(_962_), .Y(_962__bF_buf3) );
	BUFX4 BUFX4_89 ( .A(_962_), .Y(_962__bF_buf2) );
	BUFX4 BUFX4_90 ( .A(_962_), .Y(_962__bF_buf1) );
	BUFX4 BUFX4_91 ( .A(_962_), .Y(_962__bF_buf0) );
	INVX8 INVX8_1 ( .A(RDY_bF_buf8), .Y(_881_) );
	NOR2X1 NOR2X1_1 ( .A(state_5_), .B(state_4_), .Y(_882_) );
	NOR2X1 NOR2X1_2 ( .A(state_0_), .B(state_1_), .Y(_883_) );
	AND2X2 AND2X2_1 ( .A(state_2_), .B(state_3_), .Y(_884_) );
	NAND3X1 NAND3X1_1 ( .A(_882__bF_buf5), .B(_883_), .C(_884_), .Y(_885_) );
	NOR2X1 NOR2X1_3 ( .A(_881__bF_buf7), .B(_885__bF_buf4), .Y(_886_) );
	INVX4 INVX4_1 ( .A(IRHOLD_valid), .Y(_887_) );
	INVX1 INVX1_1 ( .A(DIHOLD_4_), .Y(_889_) );
	NAND2X1 NAND2X1_1 ( .A(RDY_bF_buf7), .B(DI[4]), .Y(_890_) );
	OAI21X1 OAI21X1_1 ( .A(RDY_bF_buf6), .B(_889_), .C(_890_), .Y(DIMUX_4_) );
	INVX4 INVX4_2 ( .A(DIMUX_4_), .Y(_891_) );
	INVX1 INVX1_2 ( .A(I), .Y(_892_) );
	INVX1 INVX1_3 ( .A(IRQ), .Y(_893_) );
	INVX2 INVX2_1 ( .A(NMI_edge), .Y(_894_) );
	NAND2X1 NAND2X1_2 ( .A(_893_), .B(_894_), .Y(_895_) );
	OAI21X1 OAI21X1_2 ( .A(_892_), .B(NMI_edge), .C(_895_), .Y(_896_) );
	OAI21X1 OAI21X1_3 ( .A(_887_), .B(IRHOLD_4_), .C(_896__bF_buf3), .Y(_897_) );
	AOI21X1 AOI21X1_1 ( .A(_887_), .B(_891_), .C(_897_), .Y(_898_) );
	INVX1 INVX1_4 ( .A(IRHOLD_3_), .Y(_899_) );
	INVX1 INVX1_5 ( .A(DIHOLD_3_), .Y(_900_) );
	NAND2X1 NAND2X1_3 ( .A(RDY_bF_buf5), .B(DI[3]), .Y(_901_) );
	OAI21X1 OAI21X1_4 ( .A(RDY_bF_buf4), .B(_900_), .C(_901_), .Y(DIMUX_3_) );
	NAND2X1 NAND2X1_4 ( .A(_887_), .B(DIMUX_3_), .Y(_902_) );
	OAI21X1 OAI21X1_5 ( .A(_887_), .B(_899_), .C(_902_), .Y(_903_) );
	NAND2X1 NAND2X1_5 ( .A(_896__bF_buf2), .B(_903_), .Y(_904_) );
	MUX2X1 MUX2X1_1 ( .A(DI[2]), .B(DIHOLD_2_), .S(RDY_bF_buf3), .Y(_905_) );
	NAND2X1 NAND2X1_6 ( .A(IRHOLD_valid), .B(IRHOLD_2_), .Y(_906_) );
	OAI21X1 OAI21X1_6 ( .A(IRHOLD_valid), .B(_905_), .C(_906_), .Y(_907_) );
	AND2X2 AND2X2_2 ( .A(_907_), .B(_896__bF_buf1), .Y(_908_) );
	NOR2X1 NOR2X1_4 ( .A(_908_), .B(_904_), .Y(_909_) );
	OAI21X1 OAI21X1_7 ( .A(I), .B(_893_), .C(_894_), .Y(_910_) );
	INVX1 INVX1_6 ( .A(DIHOLD_1_), .Y(_911_) );
	NAND2X1 NAND2X1_7 ( .A(RDY_bF_buf2), .B(DI[1]), .Y(_912_) );
	OAI21X1 OAI21X1_8 ( .A(RDY_bF_buf1), .B(_911_), .C(_912_), .Y(DIMUX_1_) );
	MUX2X1 MUX2X1_2 ( .A(DIMUX_1_), .B(IRHOLD_1_), .S(_887_), .Y(_913_) );
	OR2X2 OR2X2_1 ( .A(_913_), .B(_910__bF_buf4), .Y(_914_) );
	INVX1 INVX1_7 ( .A(DIHOLD_0_), .Y(_915_) );
	NAND2X1 NAND2X1_8 ( .A(RDY_bF_buf0), .B(DI[0]), .Y(_916_) );
	OAI21X1 OAI21X1_9 ( .A(RDY_bF_buf8), .B(_915_), .C(_916_), .Y(DIMUX_0_) );
	MUX2X1 MUX2X1_3 ( .A(DIMUX_0_), .B(IRHOLD_0_), .S(_887_), .Y(_917_) );
	NOR2X1 NOR2X1_5 ( .A(_910__bF_buf3), .B(_917_), .Y(_918_) );
	AND2X2 AND2X2_3 ( .A(_914_), .B(_918_), .Y(_919_) );
	NAND2X1 NAND2X1_9 ( .A(_909_), .B(_919_), .Y(_920_) );
	OAI21X1 OAI21X1_10 ( .A(_907_), .B(_903_), .C(_896__bF_buf0), .Y(_921_) );
	INVX1 INVX1_8 ( .A(IRHOLD_4_), .Y(_922_) );
	AOI21X1 AOI21X1_2 ( .A(IRHOLD_valid), .B(_922_), .C(_910__bF_buf2), .Y(_923_) );
	OAI21X1 OAI21X1_11 ( .A(IRHOLD_valid), .B(DIMUX_4_), .C(_923_), .Y(_924_) );
	MUX2X1 MUX2X1_4 ( .A(DI[7]), .B(DIHOLD_7_), .S(RDY_bF_buf7), .Y(_925_) );
	NAND2X1 NAND2X1_10 ( .A(IRHOLD_valid), .B(IRHOLD_7_), .Y(_926_) );
	OAI21X1 OAI21X1_12 ( .A(IRHOLD_valid), .B(_925_), .C(_926_), .Y(_927_) );
	AND2X2 AND2X2_4 ( .A(_927_), .B(_896__bF_buf3), .Y(_928_) );
	NAND2X1 NAND2X1_11 ( .A(_924_), .B(_928_), .Y(_929_) );
	NOR2X1 NOR2X1_6 ( .A(_918_), .B(_929_), .Y(_930_) );
	NAND2X1 NAND2X1_12 ( .A(_921_), .B(_930_), .Y(_931_) );
	OAI21X1 OAI21X1_13 ( .A(_898_), .B(_920_), .C(_931_), .Y(_932_) );
	INVX2 INVX2_2 ( .A(state_0_), .Y(_933_) );
	NOR2X1 NOR2X1_7 ( .A(state_1_), .B(_933_), .Y(_934_) );
	NOR2X1 NOR2X1_8 ( .A(state_2_), .B(state_3_), .Y(_935_) );
	NAND2X1 NAND2X1_13 ( .A(_935_), .B(_934_), .Y(_936_) );
	INVX8 INVX8_2 ( .A(_882__bF_buf4), .Y(_937_) );
	INVX1 INVX1_9 ( .A(state_3_), .Y(_938_) );
	NAND2X1 NAND2X1_14 ( .A(state_2_), .B(_938_), .Y(_939_) );
	OR2X2 OR2X2_2 ( .A(state_0_), .B(state_1_), .Y(_940_) );
	NOR2X1 NOR2X1_9 ( .A(_940_), .B(_939_), .Y(_941_) );
	NAND2X1 NAND2X1_15 ( .A(_882__bF_buf3), .B(_941_), .Y(_942_) );
	OAI21X1 OAI21X1_14 ( .A(_936__bF_buf3), .B(_937__bF_buf4), .C(_942_), .Y(_943_) );
	AND2X2 AND2X2_5 ( .A(state_5_), .B(state_4_), .Y(_944_) );
	INVX2 INVX2_3 ( .A(_944_), .Y(_945_) );
	INVX1 INVX1_10 ( .A(state_5_), .Y(_946_) );
	NOR2X1 NOR2X1_10 ( .A(state_4_), .B(_946_), .Y(_947_) );
	NAND2X1 NAND2X1_16 ( .A(state_2_), .B(state_3_), .Y(_948_) );
	NAND2X1 NAND2X1_17 ( .A(state_0_), .B(state_1_), .Y(_949_) );
	NOR2X1 NOR2X1_11 ( .A(_948_), .B(_949_), .Y(_950_) );
	NAND2X1 NAND2X1_18 ( .A(_947_), .B(_950_), .Y(_951_) );
	OAI21X1 OAI21X1_15 ( .A(_945_), .B(_936__bF_buf2), .C(_951_), .Y(_952_) );
	NOR2X1 NOR2X1_12 ( .A(_952_), .B(_943_), .Y(_953_) );
	INVX1 INVX1_11 ( .A(_936__bF_buf1), .Y(_954_) );
	INVX2 INVX2_4 ( .A(state_4_), .Y(_955_) );
	NOR2X1 NOR2X1_13 ( .A(state_5_), .B(_955_), .Y(_956_) );
	NAND2X1 NAND2X1_19 ( .A(state_5_), .B(_955_), .Y(_957_) );
	NAND3X1 NAND3X1_2 ( .A(_933_), .B(state_1_), .C(_884_), .Y(_958_) );
	NOR2X1 NOR2X1_14 ( .A(_957__bF_buf4), .B(_958_), .Y(_959_) );
	AOI21X1 AOI21X1_3 ( .A(_954_), .B(_956_), .C(_959_), .Y(_960_) );
	NOR3X1 NOR3X1_1 ( .A(state_1_), .B(_933_), .C(_948_), .Y(_961_) );
	NAND2X1 NAND2X1_20 ( .A(state_4_), .B(_946_), .Y(_962_) );
	NAND2X1 NAND2X1_21 ( .A(_957__bF_buf3), .B(_962__bF_buf4), .Y(_963_) );
	INVX2 INVX2_5 ( .A(state_2_), .Y(_964_) );
	NOR2X1 NOR2X1_15 ( .A(state_3_), .B(_964_), .Y(_965_) );
	NAND2X1 NAND2X1_22 ( .A(_934_), .B(_965_), .Y(_966_) );
	NOR2X1 NOR2X1_16 ( .A(_962__bF_buf3), .B(_966_), .Y(_967_) );
	AOI21X1 AOI21X1_4 ( .A(_961_), .B(_963_), .C(_967_), .Y(_968_) );
	NAND2X1 NAND2X1_23 ( .A(_960_), .B(_968_), .Y(_969_) );
	NAND3X1 NAND3X1_3 ( .A(RDY_bF_buf6), .B(_953_), .C(_969_), .Y(_970_) );
	NAND2X1 NAND2X1_24 ( .A(_884_), .B(_934_), .Y(_971_) );
	NOR3X1 NOR3X1_2 ( .A(state_0_), .B(state_1_), .C(_948_), .Y(_972_) );
	NAND2X1 NAND2X1_25 ( .A(RDY_bF_buf5), .B(_972_), .Y(_973_) );
	OAI21X1 OAI21X1_16 ( .A(RDY_bF_buf4), .B(_971_), .C(_973_), .Y(_974_) );
	AND2X2 AND2X2_6 ( .A(_974_), .B(_947_), .Y(_975_) );
	NAND2X1 NAND2X1_26 ( .A(_956_), .B(_941_), .Y(_976_) );
	NOR2X1 NOR2X1_17 ( .A(_937__bF_buf3), .B(_971_), .Y(_977_) );
	INVX2 INVX2_6 ( .A(_977_), .Y(_978_) );
	NOR2X1 NOR2X1_18 ( .A(ALU_CO), .B(store), .Y(_979_) );
	NAND2X1 NAND2X1_27 ( .A(RDY_bF_buf3), .B(_979_), .Y(_980_) );
	OAI22X1 OAI22X1_1 ( .A(_976_), .B(_980_), .C(RDY_bF_buf2), .D(_978_), .Y(_981_) );
	AND2X2 AND2X2_7 ( .A(state_0_), .B(state_1_), .Y(_982_) );
	NAND2X1 NAND2X1_28 ( .A(_935_), .B(_982_), .Y(_983_) );
	INVX1 INVX1_12 ( .A(_983_), .Y(_984_) );
	NAND2X1 NAND2X1_29 ( .A(_882__bF_buf2), .B(_984_), .Y(_985_) );
	INVX2 INVX2_7 ( .A(write_back), .Y(_986_) );
	NAND3X1 NAND3X1_4 ( .A(_986_), .B(RDY_bF_buf1), .C(_979_), .Y(_987_) );
	NOR2X1 NOR2X1_19 ( .A(_987_), .B(_985_), .Y(_988_) );
	NOR3X1 NOR3X1_3 ( .A(_988_), .B(_975_), .C(_981_), .Y(_989_) );
	OR2X2 OR2X2_3 ( .A(_943_), .B(_952_), .Y(_990_) );
	NAND3X1 NAND3X1_5 ( .A(_986_), .B(RDY_bF_buf0), .C(_990_), .Y(_991_) );
	NAND3X1 NAND3X1_6 ( .A(_970_), .B(_991_), .C(_989_), .Y(_992_) );
	AOI21X1 AOI21X1_5 ( .A(_932_), .B(_886__bF_buf4), .C(_992_), .Y(_993_) );
	NOR2X1 NOR2X1_20 ( .A(_910__bF_buf1), .B(_913_), .Y(_994_) );
	NOR2X1 NOR2X1_21 ( .A(_994_), .B(_918_), .Y(_995_) );
	NAND2X1 NAND2X1_30 ( .A(_921_), .B(_995_), .Y(_996_) );
	NAND2X1 NAND2X1_31 ( .A(_887_), .B(DIMUX_4_), .Y(_997_) );
	OAI21X1 OAI21X1_17 ( .A(_887_), .B(_922_), .C(_997_), .Y(_998_) );
	OAI21X1 OAI21X1_18 ( .A(_927_), .B(_998_), .C(_896__bF_buf2), .Y(_999_) );
	INVX1 INVX1_13 ( .A(DIHOLD_5_), .Y(_1000_) );
	NAND2X1 NAND2X1_32 ( .A(RDY_bF_buf8), .B(DI[5]), .Y(_1001_) );
	OAI21X1 OAI21X1_19 ( .A(RDY_bF_buf7), .B(_1000_), .C(_1001_), .Y(DIMUX_5_) );
	MUX2X1 MUX2X1_5 ( .A(DIMUX_5_), .B(IRHOLD_5_), .S(_887_), .Y(_1002_) );
	NOR2X1 NOR2X1_22 ( .A(_910__bF_buf0), .B(_1002_), .Y(_1003_) );
	INVX1 INVX1_14 ( .A(DIHOLD_6_), .Y(_1004_) );
	NAND2X1 NAND2X1_33 ( .A(RDY_bF_buf6), .B(DI[6]), .Y(_1005_) );
	OAI21X1 OAI21X1_20 ( .A(RDY_bF_buf5), .B(_1004_), .C(_1005_), .Y(DIMUX_6_) );
	INVX1 INVX1_15 ( .A(IRHOLD_6_), .Y(_1006_) );
	AOI21X1 AOI21X1_6 ( .A(IRHOLD_valid), .B(_1006_), .C(_910__bF_buf4), .Y(_1007_) );
	OAI21X1 OAI21X1_21 ( .A(IRHOLD_valid), .B(DIMUX_6_), .C(_1007_), .Y(_1008_) );
	NOR2X1 NOR2X1_23 ( .A(_1008_), .B(_1003_), .Y(_1009_) );
	NAND2X1 NAND2X1_34 ( .A(_999_), .B(_1009_), .Y(_1010_) );
	NOR2X1 NOR2X1_24 ( .A(_1010_), .B(_996_), .Y(_1011_) );
	NAND3X1 NAND3X1_7 ( .A(_934_), .B(_947_), .C(_965_), .Y(_1012_) );
	INVX1 INVX1_16 ( .A(_1012_), .Y(_1013_) );
	AOI22X1 AOI22X1_1 ( .A(_881__bF_buf6), .B(_1013_), .C(_886__bF_buf3), .D(_1011_), .Y(_1014_) );
	NAND2X1 NAND2X1_35 ( .A(_881__bF_buf5), .B(_967_), .Y(_1015_) );
	OAI21X1 OAI21X1_22 ( .A(ALU_CO), .B(store), .C(RDY_bF_buf4), .Y(_1016_) );
	OAI21X1 OAI21X1_23 ( .A(_976_), .B(_1016_), .C(_1015_), .Y(_1017_) );
	INVX1 INVX1_17 ( .A(_1017_), .Y(_1018_) );
	NAND3X1 NAND3X1_8 ( .A(_1014_), .B(_1018_), .C(_993_), .Y(_1019_) );
	INVX1 INVX1_18 ( .A(_951_), .Y(_1020_) );
	OAI21X1 OAI21X1_24 ( .A(_998_), .B(_903_), .C(_896__bF_buf1), .Y(_1021_) );
	INVX8 INVX8_3 ( .A(_886__bF_buf2), .Y(_1022_) );
	NAND2X1 NAND2X1_36 ( .A(_896__bF_buf0), .B(_907_), .Y(_1023_) );
	NOR2X1 NOR2X1_25 ( .A(_1023_), .B(_1022__bF_buf3), .Y(_1024_) );
	AOI22X1 AOI22X1_2 ( .A(_881__bF_buf4), .B(_1020_), .C(_1021_), .D(_1024_), .Y(_1025_) );
	OAI21X1 OAI21X1_25 ( .A(_937__bF_buf2), .B(_958_), .C(RDY_bF_buf3), .Y(_1026_) );
	NAND2X1 NAND2X1_37 ( .A(_884_), .B(_982_), .Y(_1027_) );
	NOR2X1 NOR2X1_26 ( .A(_937__bF_buf1), .B(_1027_), .Y(_1028_) );
	OAI21X1 OAI21X1_26 ( .A(RDY_bF_buf2), .B(_1028_), .C(_1026_), .Y(_1029_) );
	NAND2X1 NAND2X1_38 ( .A(_1029_), .B(_1025_), .Y(_1030_) );
	NAND2X1 NAND2X1_39 ( .A(_982_), .B(_965_), .Y(_1031_) );
	NOR2X1 NOR2X1_27 ( .A(_962__bF_buf2), .B(_1031_), .Y(_1032_) );
	NAND2X1 NAND2X1_40 ( .A(state_1_), .B(_933_), .Y(_1033_) );
	NOR2X1 NOR2X1_28 ( .A(_939_), .B(_1033_), .Y(_1034_) );
	INVX1 INVX1_19 ( .A(_1034__bF_buf3), .Y(_1035_) );
	OAI21X1 OAI21X1_27 ( .A(_962__bF_buf1), .B(_1035_), .C(RDY_bF_buf1), .Y(_1036_) );
	OAI21X1 OAI21X1_28 ( .A(RDY_bF_buf0), .B(_1032_), .C(_1036_), .Y(_1037_) );
	NOR2X1 NOR2X1_29 ( .A(_957__bF_buf2), .B(_1031_), .Y(_1038_) );
	OAI21X1 OAI21X1_29 ( .A(_957__bF_buf1), .B(_1035_), .C(RDY_bF_buf8), .Y(_1039_) );
	OAI21X1 OAI21X1_30 ( .A(RDY_bF_buf7), .B(_1038_), .C(_1039_), .Y(_1040_) );
	NAND2X1 NAND2X1_41 ( .A(_1037_), .B(_1040_), .Y(_1041_) );
	NOR2X1 NOR2X1_30 ( .A(_1041_), .B(_1030_), .Y(_1042_) );
	NOR3X1 NOR3X1_4 ( .A(state_2_), .B(_938_), .C(_949_), .Y(_1043_) );
	NAND2X1 NAND2X1_42 ( .A(_947_), .B(_1043_), .Y(_1044_) );
	NAND2X1 NAND2X1_43 ( .A(state_3_), .B(_964_), .Y(_1045_) );
	NOR2X1 NOR2X1_31 ( .A(_1033_), .B(_1045_), .Y(_1046_) );
	NAND2X1 NAND2X1_44 ( .A(_947_), .B(_1046_), .Y(_1047_) );
	INVX1 INVX1_20 ( .A(_1047_), .Y(_1048_) );
	NAND2X1 NAND2X1_45 ( .A(RDY_bF_buf6), .B(_1048_), .Y(_1049_) );
	OAI21X1 OAI21X1_31 ( .A(RDY_bF_buf5), .B(_1044_), .C(_1049_), .Y(_1050_) );
	NAND3X1 NAND3X1_9 ( .A(_964_), .B(state_3_), .C(_982_), .Y(_1051_) );
	NOR2X1 NOR2X1_32 ( .A(_937__bF_buf0), .B(_1051_), .Y(_1052_) );
	INVX1 INVX1_21 ( .A(_1052_), .Y(_1053_) );
	INVX1 INVX1_22 ( .A(state_1_), .Y(_1054_) );
	NOR2X1 NOR2X1_33 ( .A(state_0_), .B(_1054_), .Y(_1055_) );
	NOR2X1 NOR2X1_34 ( .A(state_2_), .B(_938_), .Y(_1056_) );
	NAND3X1 NAND3X1_10 ( .A(_882__bF_buf1), .B(_1055_), .C(_1056_), .Y(_1057_) );
	MUX2X1 MUX2X1_6 ( .A(_1053_), .B(_1057__bF_buf3), .S(_881__bF_buf3), .Y(_1058_) );
	NOR2X1 NOR2X1_35 ( .A(_1058_), .B(_1050_), .Y(_1059_) );
	OAI21X1 OAI21X1_32 ( .A(_962__bF_buf0), .B(_1051_), .C(_881__bF_buf2), .Y(_1060_) );
	NAND2X1 NAND2X1_46 ( .A(_1055_), .B(_1056_), .Y(_1061_) );
	NOR2X1 NOR2X1_36 ( .A(_962__bF_buf4), .B(_1061_), .Y(_1062_) );
	OAI21X1 OAI21X1_33 ( .A(_881__bF_buf1), .B(_1062_), .C(_1060_), .Y(_1063_) );
	NAND3X1 NAND3X1_11 ( .A(_882__bF_buf0), .B(_965_), .C(_1055_), .Y(_1064_) );
	XOR2X1 XOR2X1_1 ( .A(ALU_CO), .B(backwards), .Y(_1065_) );
	INVX1 INVX1_23 ( .A(_1065_), .Y(_1066_) );
	OAI21X1 OAI21X1_34 ( .A(_1064_), .B(_1066_), .C(RDY_bF_buf4), .Y(_1067_) );
	NOR2X1 NOR2X1_37 ( .A(_937__bF_buf4), .B(_1031_), .Y(_1068_) );
	OAI21X1 OAI21X1_35 ( .A(RDY_bF_buf3), .B(_1068_), .C(_1067_), .Y(_1069_) );
	AND2X2 AND2X2_8 ( .A(_1069_), .B(_1063_), .Y(_1070_) );
	AND2X2 AND2X2_9 ( .A(_1059_), .B(_1070_), .Y(_1071_) );
	NOR2X1 NOR2X1_38 ( .A(_986_), .B(_881__bF_buf0), .Y(_1072_) );
	NOR2X1 NOR2X1_39 ( .A(_957__bF_buf0), .B(_983_), .Y(_1073_) );
	AOI22X1 AOI22X1_3 ( .A(_881__bF_buf7), .B(_1073_), .C(_1072_), .D(_990_), .Y(_1074_) );
	NOR2X1 NOR2X1_40 ( .A(_962__bF_buf3), .B(_983_), .Y(_1075_) );
	NAND3X1 NAND3X1_12 ( .A(_933_), .B(state_1_), .C(_935_), .Y(_1076_) );
	OAI21X1 OAI21X1_36 ( .A(_962__bF_buf2), .B(_1076_), .C(RDY_bF_buf2), .Y(_1077_) );
	OAI21X1 OAI21X1_37 ( .A(RDY_bF_buf1), .B(_1075_), .C(_1077_), .Y(_1078_) );
	NAND2X1 NAND2X1_47 ( .A(_1078_), .B(_1074_), .Y(_1079_) );
	NAND3X1 NAND3X1_13 ( .A(_884_), .B(_956_), .C(_1055_), .Y(_1080_) );
	INVX1 INVX1_24 ( .A(_1080_), .Y(_1081_) );
	OAI21X1 OAI21X1_38 ( .A(_962__bF_buf1), .B(_1027_), .C(_881__bF_buf6), .Y(_1082_) );
	OAI21X1 OAI21X1_39 ( .A(_881__bF_buf5), .B(_1081_), .C(_1082_), .Y(_1083_) );
	OAI21X1 OAI21X1_40 ( .A(_937__bF_buf3), .B(_983_), .C(_881__bF_buf4), .Y(_1084_) );
	NOR2X1 NOR2X1_41 ( .A(_937__bF_buf2), .B(_1076_), .Y(_1085_) );
	OAI21X1 OAI21X1_41 ( .A(_881__bF_buf3), .B(_1085_), .C(_1084_), .Y(_1086_) );
	NAND2X1 NAND2X1_48 ( .A(_1086_), .B(_1083_), .Y(_1087_) );
	NOR2X1 NOR2X1_42 ( .A(_1087_), .B(_1079_), .Y(_1088_) );
	NAND3X1 NAND3X1_14 ( .A(_1042_), .B(_1071_), .C(_1088_), .Y(_1089_) );
	NOR2X1 NOR2X1_43 ( .A(_957__bF_buf4), .B(_936__bF_buf0), .Y(_1090_) );
	NAND2X1 NAND2X1_49 ( .A(_881__bF_buf2), .B(_1090_), .Y(_1091_) );
	NAND2X1 NAND2X1_50 ( .A(_896__bF_buf3), .B(_927_), .Y(_1092_) );
	NAND2X1 NAND2X1_51 ( .A(_1092_), .B(_924_), .Y(_1093_) );
	NOR2X1 NOR2X1_44 ( .A(_1003_), .B(_1093_), .Y(_1094_) );
	INVX4 INVX4_3 ( .A(DIMUX_3_), .Y(_1095_) );
	OAI21X1 OAI21X1_42 ( .A(_887_), .B(IRHOLD_3_), .C(_896__bF_buf2), .Y(_1096_) );
	AOI21X1 AOI21X1_7 ( .A(_887_), .B(_1095_), .C(_1096_), .Y(_1097_) );
	NAND2X1 NAND2X1_52 ( .A(_1023_), .B(_1097_), .Y(_1098_) );
	OAI21X1 OAI21X1_43 ( .A(_910__bF_buf3), .B(_917_), .C(_914_), .Y(_1099_) );
	NOR2X1 NOR2X1_45 ( .A(_1098_), .B(_1099_), .Y(_1100_) );
	NAND3X1 NAND3X1_15 ( .A(_886__bF_buf1), .B(_1094_), .C(_1100_), .Y(_1101_) );
	AND2X2 AND2X2_10 ( .A(_1101_), .B(_1091_), .Y(_1102_) );
	NAND3X1 NAND3X1_16 ( .A(_882__bF_buf5), .B(_934_), .C(_965_), .Y(_1103_) );
	INVX1 INVX1_25 ( .A(_1103_), .Y(_1104_) );
	NOR2X1 NOR2X1_46 ( .A(_924_), .B(_996_), .Y(_1105_) );
	AOI22X1 AOI22X1_4 ( .A(_881__bF_buf1), .B(_1104_), .C(_886__bF_buf0), .D(_1105_), .Y(_1106_) );
	NAND3X1 NAND3X1_17 ( .A(_935_), .B(_883_), .C(_944_), .Y(_1107_) );
	INVX1 INVX1_26 ( .A(_1107_), .Y(_1108_) );
	OAI21X1 OAI21X1_44 ( .A(_945_), .B(_936__bF_buf3), .C(_881__bF_buf0), .Y(_1109_) );
	OAI21X1 OAI21X1_45 ( .A(_881__bF_buf7), .B(_1108_), .C(_1109_), .Y(_1110_) );
	NAND2X1 NAND2X1_53 ( .A(_935_), .B(_883_), .Y(_1111_) );
	NOR2X1 NOR2X1_47 ( .A(_962__bF_buf0), .B(_1111_), .Y(_1112_) );
	OAI21X1 OAI21X1_46 ( .A(_962__bF_buf4), .B(_936__bF_buf2), .C(_881__bF_buf6), .Y(_1113_) );
	OAI21X1 OAI21X1_47 ( .A(_881__bF_buf5), .B(_1112_), .C(_1113_), .Y(_1114_) );
	NAND2X1 NAND2X1_54 ( .A(_1114_), .B(_1110_), .Y(_1115_) );
	INVX1 INVX1_27 ( .A(_1115_), .Y(_1116_) );
	NAND2X1 NAND2X1_55 ( .A(_934_), .B(_1056_), .Y(_1117_) );
	OAI21X1 OAI21X1_48 ( .A(_957__bF_buf3), .B(_1117_), .C(_881__bF_buf4), .Y(_1118_) );
	NAND3X1 NAND3X1_18 ( .A(_964_), .B(state_3_), .C(_883_), .Y(_1119_) );
	NOR2X1 NOR2X1_48 ( .A(_957__bF_buf2), .B(_1119_), .Y(_1120_) );
	OAI21X1 OAI21X1_49 ( .A(_881__bF_buf3), .B(_1120_), .C(_1118_), .Y(_1121_) );
	NOR2X1 NOR2X1_49 ( .A(_937__bF_buf1), .B(_1117_), .Y(_1122_) );
	NOR2X1 NOR2X1_50 ( .A(RDY_bF_buf0), .B(_1122_), .Y(_1123_) );
	NOR2X1 NOR2X1_51 ( .A(_940_), .B(_1045_), .Y(_1124_) );
	AOI21X1 AOI21X1_8 ( .A(_1124_), .B(_882__bF_buf4), .C(_881__bF_buf2), .Y(_1125_) );
	OAI21X1 OAI21X1_50 ( .A(_1125_), .B(_1123_), .C(_1121_), .Y(_1126_) );
	NAND3X1 NAND3X1_19 ( .A(_935_), .B(_882__bF_buf3), .C(_883_), .Y(_1127_) );
	INVX1 INVX1_28 ( .A(_1127_), .Y(_1128_) );
	OAI21X1 OAI21X1_51 ( .A(_937__bF_buf0), .B(_936__bF_buf1), .C(_881__bF_buf1), .Y(_1129_) );
	OAI21X1 OAI21X1_52 ( .A(_881__bF_buf0), .B(_1128_), .C(_1129_), .Y(_1130_) );
	OAI21X1 OAI21X1_53 ( .A(_962__bF_buf3), .B(_1117_), .C(_881__bF_buf7), .Y(_1131_) );
	NOR2X1 NOR2X1_52 ( .A(_962__bF_buf2), .B(_1119_), .Y(_1132_) );
	OAI21X1 OAI21X1_54 ( .A(_881__bF_buf6), .B(_1132_), .C(_1131_), .Y(_1133_) );
	NAND2X1 NAND2X1_56 ( .A(_956_), .B(_974_), .Y(_1134_) );
	NAND3X1 NAND3X1_20 ( .A(_1130_), .B(_1133_), .C(_1134_), .Y(_1135_) );
	NOR2X1 NOR2X1_53 ( .A(_1135_), .B(_1126_), .Y(_1136_) );
	AND2X2 AND2X2_11 ( .A(_1136_), .B(_1116_), .Y(_1137_) );
	NAND3X1 NAND3X1_21 ( .A(_1106_), .B(_1137_), .C(_1102_), .Y(_1138_) );
	NOR3X1 NOR3X1_5 ( .A(_1138_), .B(_1089_), .C(_1019_), .Y(_1139_) );
	INVX1 INVX1_29 ( .A(_1139_), .Y(_876_) );
	INVX1 INVX1_30 ( .A(_1089_), .Y(_1140_) );
	NAND2X1 NAND2X1_57 ( .A(_924_), .B(_1003_), .Y(_1141_) );
	NOR2X1 NOR2X1_54 ( .A(_928_), .B(_1141_), .Y(_1142_) );
	NAND3X1 NAND3X1_22 ( .A(_886__bF_buf4), .B(_1142_), .C(_1100_), .Y(_1143_) );
	NAND2X1 NAND2X1_58 ( .A(_881__bF_buf5), .B(_1081_), .Y(_1144_) );
	OAI21X1 OAI21X1_55 ( .A(_957__bF_buf1), .B(_958_), .C(_881__bF_buf4), .Y(_1145_) );
	OAI21X1 OAI21X1_56 ( .A(_881__bF_buf3), .B(_1073_), .C(_1145_), .Y(_1146_) );
	NAND3X1 NAND3X1_23 ( .A(_1144_), .B(_1146_), .C(_1143_), .Y(_1147_) );
	NOR2X1 NOR2X1_55 ( .A(_1023_), .B(_918_), .Y(_1148_) );
	NAND3X1 NAND3X1_24 ( .A(_1097_), .B(_914_), .C(_1148_), .Y(_1149_) );
	NOR2X1 NOR2X1_56 ( .A(_1010_), .B(_1149_), .Y(_1150_) );
	NAND2X1 NAND2X1_59 ( .A(_956_), .B(_1034__bF_buf2), .Y(_1151_) );
	NOR2X1 NOR2X1_57 ( .A(_962__bF_buf1), .B(_1117_), .Y(_1152_) );
	OAI21X1 OAI21X1_57 ( .A(_1052_), .B(_1152_), .C(RDY_bF_buf8), .Y(_1153_) );
	OAI21X1 OAI21X1_58 ( .A(RDY_bF_buf7), .B(_1151_), .C(_1153_), .Y(_1154_) );
	AOI21X1 AOI21X1_9 ( .A(_1150_), .B(_886__bF_buf3), .C(_1154_), .Y(_1155_) );
	NOR2X1 NOR2X1_58 ( .A(_937__bF_buf4), .B(_958_), .Y(_1156_) );
	NAND2X1 NAND2X1_60 ( .A(_881__bF_buf2), .B(_1156_), .Y(_1157_) );
	NAND2X1 NAND2X1_61 ( .A(_921_), .B(_919_), .Y(_1158_) );
	NOR2X1 NOR2X1_59 ( .A(_898_), .B(_1158_), .Y(_1159_) );
	NAND2X1 NAND2X1_62 ( .A(_886__bF_buf2), .B(_1159_), .Y(_1160_) );
	NAND3X1 NAND3X1_25 ( .A(_1157_), .B(_1160_), .C(_1155_), .Y(_1161_) );
	OR2X2 OR2X2_4 ( .A(_1002_), .B(_910__bF_buf2), .Y(_1162_) );
	NOR2X1 NOR2X1_60 ( .A(_898_), .B(_1162_), .Y(_1163_) );
	NAND2X1 NAND2X1_63 ( .A(_1092_), .B(_1008_), .Y(_1164_) );
	INVX1 INVX1_31 ( .A(_1164_), .Y(_1165_) );
	NAND2X1 NAND2X1_64 ( .A(_1165_), .B(_1163_), .Y(_1166_) );
	NOR2X1 NOR2X1_61 ( .A(_996_), .B(_1166_), .Y(_1167_) );
	AOI22X1 AOI22X1_5 ( .A(_881__bF_buf1), .B(_1062_), .C(_886__bF_buf1), .D(_1167_), .Y(_1168_) );
	NOR2X1 NOR2X1_62 ( .A(_1008_), .B(_928_), .Y(_1169_) );
	NAND2X1 NAND2X1_65 ( .A(_1169_), .B(_1163_), .Y(_1170_) );
	NOR2X1 NOR2X1_63 ( .A(_996_), .B(_1170_), .Y(_1171_) );
	AOI22X1 AOI22X1_6 ( .A(_881__bF_buf0), .B(_1048_), .C(_886__bF_buf0), .D(_1171_), .Y(_1172_) );
	NOR2X1 NOR2X1_64 ( .A(_881__bF_buf7), .B(_1103_), .Y(_1173_) );
	INVX1 INVX1_32 ( .A(Z), .Y(_1174_) );
	NAND2X1 NAND2X1_66 ( .A(cond_code_1_), .B(_1174_), .Y(_1175_) );
	OAI21X1 OAI21X1_59 ( .A(cond_code_1_), .B(C), .C(_1175_), .Y(_1176_) );
	INVX1 INVX1_33 ( .A(V), .Y(_1177_) );
	NAND2X1 NAND2X1_67 ( .A(cond_code_1_), .B(_1177_), .Y(_1178_) );
	OAI21X1 OAI21X1_60 ( .A(N), .B(cond_code_1_), .C(_1178_), .Y(_1179_) );
	MUX2X1 MUX2X1_7 ( .A(_1176_), .B(_1179_), .S(cond_code_2_), .Y(_1180_) );
	XNOR2X1 XNOR2X1_1 ( .A(_1180_), .B(cond_code_0_), .Y(_1181_) );
	OAI21X1 OAI21X1_61 ( .A(_957__bF_buf0), .B(_1035_), .C(_881__bF_buf6), .Y(_1182_) );
	OAI21X1 OAI21X1_62 ( .A(_881__bF_buf5), .B(_1013_), .C(_1182_), .Y(_1183_) );
	OAI21X1 OAI21X1_63 ( .A(RDY_bF_buf6), .B(_1064_), .C(_1183_), .Y(_1184_) );
	AOI21X1 AOI21X1_10 ( .A(_1181_), .B(_1173_), .C(_1184_), .Y(_1185_) );
	NAND3X1 NAND3X1_26 ( .A(_1185_), .B(_1168_), .C(_1172_), .Y(_1186_) );
	NOR3X1 NOR3X1_6 ( .A(_1147_), .B(_1161_), .C(_1186_), .Y(_1187_) );
	NOR2X1 NOR2X1_65 ( .A(_962__bF_buf0), .B(_1076_), .Y(_1188_) );
	NOR2X1 NOR2X1_66 ( .A(_924_), .B(_1158_), .Y(_1189_) );
	AOI22X1 AOI22X1_7 ( .A(_881__bF_buf4), .B(_1188_), .C(_886__bF_buf4), .D(_1189_), .Y(_1190_) );
	NAND2X1 NAND2X1_68 ( .A(state_0_), .B(_1054_), .Y(_1191_) );
	NOR2X1 NOR2X1_67 ( .A(_1191_), .B(_1045_), .Y(_1192_) );
	NAND2X1 NAND2X1_69 ( .A(_882__bF_buf2), .B(_1192_), .Y(_1193_) );
	INVX2 INVX2_8 ( .A(_1057__bF_buf2), .Y(_1194_) );
	NAND2X1 NAND2X1_70 ( .A(_881__bF_buf3), .B(_1194_), .Y(_1195_) );
	OAI21X1 OAI21X1_64 ( .A(_881__bF_buf2), .B(_1193_), .C(_1195_), .Y(_1196_) );
	INVX1 INVX1_34 ( .A(_1085_), .Y(_1197_) );
	NOR2X1 NOR2X1_68 ( .A(_957__bF_buf4), .B(_1076_), .Y(_1198_) );
	OAI21X1 OAI21X1_65 ( .A(_957__bF_buf3), .B(_936__bF_buf0), .C(RDY_bF_buf5), .Y(_1199_) );
	OAI21X1 OAI21X1_66 ( .A(RDY_bF_buf4), .B(_1198_), .C(_1199_), .Y(_1200_) );
	OAI21X1 OAI21X1_67 ( .A(RDY_bF_buf3), .B(_1197_), .C(_1200_), .Y(_1201_) );
	OR2X2 OR2X2_5 ( .A(_1201_), .B(_1196_), .Y(_1202_) );
	OAI21X1 OAI21X1_68 ( .A(_910__bF_buf1), .B(_913_), .C(_918_), .Y(_1203_) );
	NAND2X1 NAND2X1_71 ( .A(_908_), .B(_1097_), .Y(_1204_) );
	OAI21X1 OAI21X1_69 ( .A(_1203_), .B(_1098_), .C(_1204_), .Y(_1205_) );
	NOR2X1 NOR2X1_69 ( .A(_924_), .B(_1022__bF_buf2), .Y(_1206_) );
	AOI21X1 AOI21X1_11 ( .A(_1205_), .B(_1206_), .C(_1202_), .Y(_1207_) );
	AND2X2 AND2X2_12 ( .A(_1190_), .B(_1207_), .Y(_1208_) );
	NAND3X1 NAND3X1_27 ( .A(_1140_), .B(_1208_), .C(_1187_), .Y(_877_) );
	NAND2X1 NAND2X1_72 ( .A(_883_), .B(_965_), .Y(_1209_) );
	OAI21X1 OAI21X1_70 ( .A(_962__bF_buf4), .B(_1209_), .C(_881__bF_buf1), .Y(_1210_) );
	OAI21X1 OAI21X1_71 ( .A(_881__bF_buf0), .B(_1075_), .C(_1210_), .Y(_1211_) );
	NOR2X1 NOR2X1_70 ( .A(_881__bF_buf7), .B(_990_), .Y(_1212_) );
	OR2X2 OR2X2_6 ( .A(state_2_), .B(state_3_), .Y(_1213_) );
	NOR2X1 NOR2X1_71 ( .A(_1213_), .B(_1033_), .Y(_1215_) );
	OAI21X1 OAI21X1_72 ( .A(_1215_), .B(_1192_), .C(_947_), .Y(_1216_) );
	OAI21X1 OAI21X1_73 ( .A(state_5_), .B(_1031_), .C(_1216_), .Y(_1217_) );
	NOR2X1 NOR2X1_72 ( .A(_957__bF_buf2), .B(_1111_), .Y(_1218_) );
	NOR2X1 NOR2X1_73 ( .A(_957__bF_buf1), .B(_1209_), .Y(_1219_) );
	NOR2X1 NOR2X1_74 ( .A(_1218_), .B(_1219_), .Y(_1220_) );
	OAI21X1 OAI21X1_74 ( .A(_937__bF_buf3), .B(_971_), .C(_1220_), .Y(_1221_) );
	OAI21X1 OAI21X1_75 ( .A(_1217_), .B(_1221_), .C(_1212_), .Y(_1222_) );
	INVX1 INVX1_35 ( .A(_1181_), .Y(_1223_) );
	INVX8 INVX8_4 ( .A(_1064_), .Y(_1224_) );
	NAND3X1 NAND3X1_28 ( .A(RDY_bF_buf2), .B(_1066_), .C(_1224_), .Y(_1225_) );
	OAI21X1 OAI21X1_76 ( .A(RDY_bF_buf1), .B(_885__bF_buf3), .C(_1225_), .Y(_1226_) );
	AOI21X1 AOI21X1_12 ( .A(_1223_), .B(_1173_), .C(_1226_), .Y(_1227_) );
	AND2X2 AND2X2_13 ( .A(_1222_), .B(_1227_), .Y(_1228_) );
	AOI21X1 AOI21X1_13 ( .A(_1010_), .B(_924_), .C(_996_), .Y(_1229_) );
	NAND2X1 NAND2X1_73 ( .A(_1094_), .B(_1100_), .Y(_1230_) );
	OAI21X1 OAI21X1_77 ( .A(_924_), .B(_1158_), .C(_1230_), .Y(_1231_) );
	NOR2X1 NOR2X1_75 ( .A(_1229_), .B(_1231_), .Y(_1232_) );
	NAND2X1 NAND2X1_74 ( .A(_1142_), .B(_1100_), .Y(_1233_) );
	OAI21X1 OAI21X1_78 ( .A(_996_), .B(_1170_), .C(_1233_), .Y(_1234_) );
	NAND2X1 NAND2X1_75 ( .A(_1023_), .B(_904_), .Y(_1235_) );
	NOR2X1 NOR2X1_76 ( .A(_1203_), .B(_1235_), .Y(_1236_) );
	NAND2X1 NAND2X1_76 ( .A(_924_), .B(_1236_), .Y(_1237_) );
	OAI21X1 OAI21X1_79 ( .A(_1149_), .B(_1170_), .C(_1237_), .Y(_1238_) );
	NOR2X1 NOR2X1_77 ( .A(_1238_), .B(_1234_), .Y(_1239_) );
	NOR2X1 NOR2X1_78 ( .A(_1203_), .B(_1098_), .Y(_1240_) );
	AOI22X1 AOI22X1_8 ( .A(_921_), .B(_930_), .C(_924_), .D(_1240_), .Y(_1241_) );
	OAI21X1 OAI21X1_80 ( .A(_1023_), .B(_1097_), .C(_886__bF_buf3), .Y(_1242_) );
	INVX1 INVX1_36 ( .A(_1242_), .Y(_1243_) );
	NAND2X1 NAND2X1_77 ( .A(_1243_), .B(_1241_), .Y(_1244_) );
	AOI21X1 AOI21X1_14 ( .A(_898_), .B(_1205_), .C(_1244_), .Y(_1245_) );
	NAND3X1 NAND3X1_29 ( .A(_1232_), .B(_1239_), .C(_1245_), .Y(_1246_) );
	NOR2X1 NOR2X1_79 ( .A(_1204_), .B(_1099_), .Y(_1247_) );
	OAI21X1 OAI21X1_81 ( .A(_1164_), .B(_1141_), .C(_929_), .Y(_1248_) );
	OAI21X1 OAI21X1_82 ( .A(_910__bF_buf0), .B(_917_), .C(_994_), .Y(_1249_) );
	NAND2X1 NAND2X1_78 ( .A(_1203_), .B(_1249_), .Y(_1250_) );
	NOR2X1 NOR2X1_80 ( .A(_898_), .B(_1204_), .Y(_1251_) );
	AND2X2 AND2X2_14 ( .A(_1251_), .B(_1250_), .Y(_1252_) );
	AOI21X1 AOI21X1_15 ( .A(_1247_), .B(_1248_), .C(_1252_), .Y(_1253_) );
	NOR2X1 NOR2X1_81 ( .A(_1249_), .B(_1098_), .Y(_1254_) );
	AOI21X1 AOI21X1_16 ( .A(_1100_), .B(_1093_), .C(_1254_), .Y(_1255_) );
	OAI21X1 OAI21X1_83 ( .A(_910__bF_buf4), .B(_1002_), .C(_924_), .Y(_1256_) );
	INVX1 INVX1_37 ( .A(_1256_), .Y(_1257_) );
	NAND2X1 NAND2X1_79 ( .A(_1165_), .B(_1257_), .Y(_1258_) );
	NOR2X1 NOR2X1_82 ( .A(_996_), .B(_1258_), .Y(_1259_) );
	INVX2 INVX2_9 ( .A(DIMUX_6_), .Y(_1260_) );
	OAI21X1 OAI21X1_84 ( .A(_887_), .B(IRHOLD_6_), .C(_896__bF_buf1), .Y(_1261_) );
	AOI21X1 AOI21X1_17 ( .A(_887_), .B(_1260_), .C(_1261_), .Y(_1262_) );
	NAND2X1 NAND2X1_80 ( .A(_1092_), .B(_1262_), .Y(_1263_) );
	NOR2X1 NOR2X1_83 ( .A(_1256_), .B(_1263_), .Y(_1264_) );
	NAND2X1 NAND2X1_81 ( .A(_1264_), .B(_1247_), .Y(_1265_) );
	OAI21X1 OAI21X1_85 ( .A(_996_), .B(_1166_), .C(_1265_), .Y(_1266_) );
	NOR2X1 NOR2X1_84 ( .A(_1259_), .B(_1266_), .Y(_1267_) );
	NAND3X1 NAND3X1_30 ( .A(_1253_), .B(_1255_), .C(_1267_), .Y(_1268_) );
	OAI21X1 OAI21X1_86 ( .A(_1268_), .B(_1246_), .C(_1228_), .Y(_1269_) );
	NAND2X1 NAND2X1_82 ( .A(_883_), .B(_884_), .Y(_1270_) );
	NOR2X1 NOR2X1_85 ( .A(_957__bF_buf0), .B(_1270_), .Y(_1271_) );
	OAI21X1 OAI21X1_87 ( .A(_957__bF_buf4), .B(_1051_), .C(RDY_bF_buf0), .Y(_1272_) );
	OAI21X1 OAI21X1_88 ( .A(RDY_bF_buf8), .B(_1271_), .C(_1272_), .Y(_1273_) );
	NOR2X1 NOR2X1_86 ( .A(_962__bF_buf3), .B(_1270_), .Y(_1274_) );
	OAI21X1 OAI21X1_89 ( .A(_962__bF_buf2), .B(_1051_), .C(RDY_bF_buf7), .Y(_1275_) );
	OAI21X1 OAI21X1_90 ( .A(RDY_bF_buf6), .B(_1274_), .C(_1275_), .Y(_1276_) );
	NAND2X1 NAND2X1_83 ( .A(_1276_), .B(_1273_), .Y(_1277_) );
	NOR2X1 NOR2X1_87 ( .A(_1277_), .B(_1269_), .Y(_1278_) );
	OR2X2 OR2X2_7 ( .A(_1161_), .B(_1147_), .Y(_1279_) );
	NAND2X1 NAND2X1_84 ( .A(_881__bF_buf6), .B(_1219_), .Y(_1280_) );
	OAI21X1 OAI21X1_91 ( .A(_1022__bF_buf1), .B(_1255_), .C(_1280_), .Y(_1281_) );
	INVX1 INVX1_38 ( .A(_942_), .Y(_1282_) );
	NAND2X1 NAND2X1_85 ( .A(write_back), .B(RDY_bF_buf5), .Y(_1283_) );
	AOI21X1 AOI21X1_18 ( .A(_1016_), .B(_1283_), .C(_985_), .Y(_1284_) );
	AOI21X1 AOI21X1_19 ( .A(_1282_), .B(_881__bF_buf5), .C(_1284_), .Y(_1285_) );
	INVX1 INVX1_39 ( .A(_1285_), .Y(_1286_) );
	NOR2X1 NOR2X1_88 ( .A(_1286_), .B(_1281_), .Y(_1287_) );
	AND2X2 AND2X2_15 ( .A(_1069_), .B(_1134_), .Y(_1288_) );
	AND2X2 AND2X2_16 ( .A(_1288_), .B(_1083_), .Y(_1289_) );
	AND2X2 AND2X2_17 ( .A(_1289_), .B(_1185_), .Y(_1290_) );
	AND2X2 AND2X2_18 ( .A(_1290_), .B(_1106_), .Y(_1291_) );
	NAND3X1 NAND3X1_31 ( .A(_1042_), .B(_1291_), .C(_1287_), .Y(_1292_) );
	NOR3X1 NOR3X1_7 ( .A(_1019_), .B(_1279_), .C(_1292_), .Y(_1293_) );
	NAND3X1 NAND3X1_32 ( .A(_1211_), .B(_1293_), .C(_1278_), .Y(_878_) );
	AOI22X1 AOI22X1_9 ( .A(_1100_), .B(_1142_), .C(_898_), .D(_1205_), .Y(_1294_) );
	NAND3X1 NAND3X1_33 ( .A(_1241_), .B(_1255_), .C(_1294_), .Y(_1295_) );
	INVX1 INVX1_40 ( .A(_1295_), .Y(_1296_) );
	NOR2X1 NOR2X1_89 ( .A(_1235_), .B(_1099_), .Y(_1297_) );
	NOR2X1 NOR2X1_90 ( .A(_1141_), .B(_1263_), .Y(_1298_) );
	NAND2X1 NAND2X1_86 ( .A(_1298_), .B(_1297_), .Y(_1299_) );
	NAND3X1 NAND3X1_34 ( .A(_1237_), .B(_1265_), .C(_1299_), .Y(_1300_) );
	INVX1 INVX1_41 ( .A(_1229_), .Y(_1301_) );
	AOI21X1 AOI21X1_20 ( .A(_1100_), .B(_1094_), .C(_1242_), .Y(_1302_) );
	NAND2X1 NAND2X1_87 ( .A(_1302_), .B(_1301_), .Y(_1303_) );
	NOR3X1 NOR3X1_8 ( .A(_1167_), .B(_1300_), .C(_1303_), .Y(_1304_) );
	NAND2X1 NAND2X1_88 ( .A(_1298_), .B(_1247_), .Y(_1305_) );
	NOR2X1 NOR2X1_91 ( .A(_1259_), .B(_1189_), .Y(_1306_) );
	NAND3X1 NAND3X1_35 ( .A(_1305_), .B(_1253_), .C(_1306_), .Y(_1307_) );
	INVX1 INVX1_42 ( .A(_1307_), .Y(_1308_) );
	NAND3X1 NAND3X1_36 ( .A(_1296_), .B(_1304_), .C(_1308_), .Y(_1309_) );
	INVX1 INVX1_43 ( .A(_1211_), .Y(_1310_) );
	NOR2X1 NOR2X1_92 ( .A(_1277_), .B(_1310_), .Y(_1311_) );
	NAND3X1 NAND3X1_37 ( .A(_1228_), .B(_1311_), .C(_1309_), .Y(_1312_) );
	NAND2X1 NAND2X1_89 ( .A(_995_), .B(_909_), .Y(_1313_) );
	NOR2X1 NOR2X1_93 ( .A(_999_), .B(_1313_), .Y(_1314_) );
	OAI21X1 OAI21X1_92 ( .A(_1254_), .B(_1314_), .C(_886__bF_buf2), .Y(_1315_) );
	NAND3X1 NAND3X1_38 ( .A(_1280_), .B(_1285_), .C(_1315_), .Y(_1316_) );
	NOR2X1 NOR2X1_94 ( .A(_1023_), .B(_1097_), .Y(_1317_) );
	AOI22X1 AOI22X1_10 ( .A(_881__bF_buf4), .B(_1108_), .C(_1206_), .D(_1317_), .Y(_1318_) );
	OAI21X1 OAI21X1_93 ( .A(_937__bF_buf2), .B(_1027_), .C(RDY_bF_buf4), .Y(_1319_) );
	OAI21X1 OAI21X1_94 ( .A(RDY_bF_buf3), .B(_1112_), .C(_1319_), .Y(_1320_) );
	NAND2X1 NAND2X1_90 ( .A(_1320_), .B(_1318_), .Y(_1321_) );
	OAI21X1 OAI21X1_95 ( .A(_962__bF_buf1), .B(_1027_), .C(RDY_bF_buf2), .Y(_1322_) );
	OAI21X1 OAI21X1_96 ( .A(RDY_bF_buf1), .B(_1218_), .C(_1322_), .Y(_1323_) );
	OAI21X1 OAI21X1_97 ( .A(RDY_bF_buf0), .B(_1127_), .C(_1323_), .Y(_1324_) );
	NOR2X1 NOR2X1_95 ( .A(_1324_), .B(_1321_), .Y(_1325_) );
	NAND3X1 NAND3X1_39 ( .A(_1207_), .B(_1325_), .C(_1190_), .Y(_1326_) );
	NAND3X1 NAND3X1_40 ( .A(_886__bF_buf1), .B(_1298_), .C(_1247_), .Y(_1327_) );
	NAND2X1 NAND2X1_91 ( .A(_881__bF_buf3), .B(_1132_), .Y(_1329_) );
	AND2X2 AND2X2_19 ( .A(_1327_), .B(_1329_), .Y(_1330_) );
	OAI21X1 OAI21X1_98 ( .A(_957__bF_buf3), .B(_1031_), .C(RDY_bF_buf8), .Y(_1331_) );
	OAI21X1 OAI21X1_99 ( .A(RDY_bF_buf7), .B(_1120_), .C(_1331_), .Y(_1332_) );
	AND2X2 AND2X2_20 ( .A(_1247_), .B(_1248_), .Y(_1333_) );
	OAI21X1 OAI21X1_100 ( .A(_1252_), .B(_1333_), .C(_886__bF_buf0), .Y(_1334_) );
	NAND3X1 NAND3X1_41 ( .A(_1330_), .B(_1332_), .C(_1334_), .Y(_1335_) );
	NOR3X1 NOR3X1_9 ( .A(_1316_), .B(_1326_), .C(_1335_), .Y(_1336_) );
	NAND3X1 NAND3X1_42 ( .A(_1187_), .B(_1336_), .C(_1139_), .Y(_1337_) );
	OAI21X1 OAI21X1_101 ( .A(_1022__bF_buf0), .B(_1237_), .C(_1157_), .Y(_1338_) );
	NOR3X1 NOR3X1_10 ( .A(_1196_), .B(_1277_), .C(_1126_), .Y(_1339_) );
	NAND2X1 NAND2X1_92 ( .A(_1083_), .B(_1063_), .Y(_1340_) );
	NAND2X1 NAND2X1_93 ( .A(_1133_), .B(_1134_), .Y(_1341_) );
	NOR2X1 NOR2X1_96 ( .A(_1341_), .B(_1340_), .Y(_1342_) );
	NAND3X1 NAND3X1_43 ( .A(_1059_), .B(_1342_), .C(_1339_), .Y(_1343_) );
	NOR3X1 NOR3X1_11 ( .A(_1030_), .B(_1343_), .C(_1338_), .Y(_1344_) );
	NAND2X1 NAND2X1_94 ( .A(_1168_), .B(_1172_), .Y(_1346_) );
	NOR2X1 NOR2X1_97 ( .A(_1147_), .B(_1346_), .Y(_1347_) );
	NOR2X1 NOR2X1_98 ( .A(_1022__bF_buf3), .B(_1241_), .Y(_1348_) );
	NAND3X1 NAND3X1_44 ( .A(_1329_), .B(_1332_), .C(_1327_), .Y(_1349_) );
	NOR3X1 NOR3X1_12 ( .A(_992_), .B(_1349_), .C(_1348_), .Y(_1350_) );
	NAND3X1 NAND3X1_45 ( .A(_1344_), .B(_1350_), .C(_1347_), .Y(_1351_) );
	NOR2X1 NOR2X1_99 ( .A(_1351_), .B(_1269_), .Y(_1353_) );
	OAI21X1 OAI21X1_102 ( .A(_1312_), .B(_1337_), .C(_1353_), .Y(_879_) );
	NAND3X1 NAND3X1_46 ( .A(_1276_), .B(_1211_), .C(_1018_), .Y(_1354_) );
	NAND2X1 NAND2X1_95 ( .A(_1078_), .B(_1037_), .Y(_1355_) );
	NOR2X1 NOR2X1_100 ( .A(_1355_), .B(_1354_), .Y(_1356_) );
	NAND3X1 NAND3X1_47 ( .A(_1116_), .B(_1342_), .C(_1356_), .Y(_1357_) );
	NOR2X1 NOR2X1_101 ( .A(_1321_), .B(_1357_), .Y(_1358_) );
	NAND3X1 NAND3X1_48 ( .A(_1190_), .B(_1330_), .C(_1358_), .Y(_1360_) );
	AND2X2 AND2X2_21 ( .A(_1143_), .B(_1144_), .Y(_1361_) );
	NAND3X1 NAND3X1_49 ( .A(_1155_), .B(_1361_), .C(_1168_), .Y(_1362_) );
	OR2X2 OR2X2_8 ( .A(_1360_), .B(_1362_), .Y(_880_) );
	NAND3X1 NAND3X1_50 ( .A(_1014_), .B(_1102_), .C(_1172_), .Y(_1364_) );
	AND2X2 AND2X2_22 ( .A(_1183_), .B(_1200_), .Y(_1365_) );
	NAND3X1 NAND3X1_51 ( .A(_1146_), .B(_1365_), .C(_1074_), .Y(_1366_) );
	NOR2X1 NOR2X1_102 ( .A(_975_), .B(_1050_), .Y(_1367_) );
	NAND3X1 NAND3X1_52 ( .A(_1110_), .B(_1121_), .C(_1367_), .Y(_1368_) );
	AND2X2 AND2X2_23 ( .A(_1332_), .B(_1273_), .Y(_1369_) );
	NAND3X1 NAND3X1_53 ( .A(_1040_), .B(_1323_), .C(_1369_), .Y(_1370_) );
	OR2X2 OR2X2_9 ( .A(_1368_), .B(_1370_), .Y(_1371_) );
	NOR2X1 NOR2X1_103 ( .A(_1366_), .B(_1371_), .Y(_1372_) );
	NAND3X1 NAND3X1_54 ( .A(_1025_), .B(_1318_), .C(_1372_), .Y(_1373_) );
	NOR2X1 NOR2X1_104 ( .A(_1364_), .B(_1373_), .Y(_1374_) );
	NAND3X1 NAND3X1_55 ( .A(_1315_), .B(_1280_), .C(_1374_), .Y(_888_) );
	INVX1 INVX1_44 ( .A(C), .Y(_1376_) );
	INVX2 INVX2_10 ( .A(shift), .Y(_1377_) );
	OAI21X1 OAI21X1_103 ( .A(_941_), .B(_984_), .C(_947_), .Y(_1378_) );
	OAI21X1 OAI21X1_104 ( .A(_937__bF_buf1), .B(_971_), .C(_1378_), .Y(_1379_) );
	NOR2X1 NOR2X1_105 ( .A(load_only), .B(_978_), .Y(_1380_) );
	AOI22X1 AOI22X1_11 ( .A(rotate), .B(_1379_), .C(_1377_), .D(_1380_), .Y(_1382_) );
	INVX1 INVX1_45 ( .A(rotate), .Y(_1383_) );
	INVX2 INVX2_11 ( .A(compare), .Y(_1384_) );
	INVX1 INVX1_46 ( .A(_1378_), .Y(_1385_) );
	NAND3X1 NAND3X1_56 ( .A(_1377_), .B(inc), .C(_1385_), .Y(_1386_) );
	OAI21X1 OAI21X1_105 ( .A(_1384_), .B(_978_), .C(_1386_), .Y(_1387_) );
	INVX1 INVX1_47 ( .A(_976_), .Y(_1388_) );
	OAI21X1 OAI21X1_106 ( .A(_937__bF_buf0), .B(_983_), .C(_1064_), .Y(_1390_) );
	OAI21X1 OAI21X1_107 ( .A(_1390_), .B(_1388_), .C(ALU_CO), .Y(_1391_) );
	INVX4 INVX4_4 ( .A(_1038_), .Y(_1392_) );
	OAI21X1 OAI21X1_108 ( .A(_937__bF_buf4), .B(_1027_), .C(_1392_), .Y(_1393_) );
	OAI21X1 OAI21X1_109 ( .A(_962__bF_buf0), .B(_1076_), .C(_1044_), .Y(_1394_) );
	NOR2X1 NOR2X1_106 ( .A(_1394_), .B(_1393_), .Y(_1395_) );
	AOI21X1 AOI21X1_21 ( .A(_947_), .B(_1034__bF_buf1), .C(_1081_), .Y(_1396_) );
	OAI21X1 OAI21X1_110 ( .A(_957__bF_buf2), .B(_1061_), .C(_1012_), .Y(_1397_) );
	INVX1 INVX1_48 ( .A(_1397_), .Y(_1398_) );
	AND2X2 AND2X2_24 ( .A(_1396_), .B(_1398_), .Y(_1399_) );
	NAND3X1 NAND3X1_57 ( .A(_1391_), .B(_1395_), .C(_1399_), .Y(_1400_) );
	AOI21X1 AOI21X1_22 ( .A(_1383_), .B(_1387_), .C(_1400_), .Y(_1401_) );
	OAI21X1 OAI21X1_111 ( .A(_1376_), .B(_1382_), .C(_1401_), .Y(ALU_CI) );
	INVX4 INVX4_5 ( .A(PC_0_), .Y(_1402_) );
	INVX2 INVX2_12 ( .A(DIMUX_0_), .Y(_1403_) );
	NOR2X1 NOR2X1_107 ( .A(_1073_), .B(_1122_), .Y(_1404_) );
	NOR2X1 NOR2X1_108 ( .A(_1224_), .B(_1062_), .Y(_1405_) );
	AOI22X1 AOI22X1_12 ( .A(_956_), .B(_972_), .C(_947_), .D(_1215_), .Y(_1406_) );
	NOR2X1 NOR2X1_109 ( .A(state_4_), .B(_1061_), .Y(_1407_) );
	NAND3X1 NAND3X1_58 ( .A(_882__bF_buf1), .B(_883_), .C(_1056_), .Y(_1408_) );
	OAI21X1 OAI21X1_112 ( .A(_957__bF_buf1), .B(_1209_), .C(_1408_), .Y(_1409_) );
	NOR2X1 NOR2X1_110 ( .A(_1407_), .B(_1409_), .Y(_1410_) );
	NAND3X1 NAND3X1_59 ( .A(_1406_), .B(_1405_), .C(_1410_), .Y(_1411_) );
	AOI21X1 AOI21X1_23 ( .A(_963_), .B(_1043_), .C(_1393_), .Y(_1412_) );
	INVX1 INVX1_49 ( .A(_966_), .Y(_1413_) );
	AOI21X1 AOI21X1_24 ( .A(_955_), .B(_1413_), .C(_1090_), .Y(_1414_) );
	NAND3X1 NAND3X1_60 ( .A(_1396_), .B(_1414_), .C(_1412_), .Y(_1415_) );
	NOR2X1 NOR2X1_111 ( .A(_1411_), .B(_1415_), .Y(_1416_) );
	NAND2X1 NAND2X1_96 ( .A(_1404_), .B(_1416_), .Y(_1417_) );
	OAI22X1 OAI22X1_2 ( .A(_1402_), .B(_1103_), .C(_1403_), .D(_1417_), .Y(ALU_BI_0_) );
	INVX2 INVX2_13 ( .A(PC_1_), .Y(_1418_) );
	INVX2 INVX2_14 ( .A(DIMUX_1_), .Y(_1419_) );
	OAI22X1 OAI22X1_3 ( .A(_1418_), .B(_1103_), .C(_1419_), .D(_1417_), .Y(ALU_BI_1_) );
	INVX1 INVX1_50 ( .A(_905_), .Y(DIMUX_2_) );
	INVX2 INVX2_15 ( .A(PC_2_), .Y(_1420_) );
	OAI22X1 OAI22X1_4 ( .A(_1420_), .B(_1103_), .C(_905_), .D(_1417_), .Y(ALU_BI_2_) );
	INVX4 INVX4_6 ( .A(PC_3_), .Y(_1421_) );
	OAI22X1 OAI22X1_5 ( .A(_1421_), .B(_1103_), .C(_1095_), .D(_1417_), .Y(ALU_BI_3_) );
	INVX2 INVX2_16 ( .A(PC_4_), .Y(_1422_) );
	OAI22X1 OAI22X1_6 ( .A(_1422_), .B(_1103_), .C(_891_), .D(_1417_), .Y(ALU_BI_4_) );
	INVX2 INVX2_17 ( .A(PC_5_), .Y(_1423_) );
	INVX1 INVX1_51 ( .A(DIMUX_5_), .Y(_1424_) );
	OAI22X1 OAI22X1_7 ( .A(_1423_), .B(_1103_), .C(_1424_), .D(_1417_), .Y(ALU_BI_5_) );
	INVX2 INVX2_18 ( .A(PC_6_), .Y(_1425_) );
	OAI22X1 OAI22X1_8 ( .A(_1425_), .B(_1103_), .C(_1260_), .D(_1417_), .Y(ALU_BI_6_) );
	INVX2 INVX2_19 ( .A(_925_), .Y(DIMUX_7_) );
	INVX2 INVX2_20 ( .A(PC_7_), .Y(_1426_) );
	OAI22X1 OAI22X1_9 ( .A(_1426_), .B(_1103_), .C(_925_), .D(_1417_), .Y(ALU_BI_7_) );
	NAND2X1 NAND2X1_97 ( .A(_947_), .B(_1034__bF_buf0), .Y(_1427_) );
	NAND3X1 NAND3X1_61 ( .A(_1057__bF_buf1), .B(_1427_), .C(_1193_), .Y(_1428_) );
	INVX1 INVX1_52 ( .A(_1428_), .Y(_1429_) );
	NAND2X1 NAND2X1_98 ( .A(_1429_), .B(_1412_), .Y(_1430_) );
	OAI21X1 OAI21X1_113 ( .A(_957__bF_buf0), .B(_983_), .C(_1103_), .Y(_1431_) );
	INVX4 INVX4_7 ( .A(_1431_), .Y(_1432_) );
	NAND3X1 NAND3X1_62 ( .A(ABH_0_), .B(_882__bF_buf0), .C(_1034__bF_buf3), .Y(_1433_) );
	OAI21X1 OAI21X1_114 ( .A(_1403_), .B(_1432_), .C(_1433_), .Y(_1434_) );
	AOI21X1 AOI21X1_25 ( .A(_1430_), .B(ADD_0_), .C(_1434_), .Y(_1435_) );
	INVX4 INVX4_8 ( .A(_885__bF_buf2), .Y(_1436_) );
	OAI22X1 OAI22X1_10 ( .A(_983_), .B(_962__bF_buf4), .C(_937__bF_buf3), .D(_958_), .Y(_1437_) );
	OAI21X1 OAI21X1_115 ( .A(_937__bF_buf2), .B(_1076_), .C(_1107_), .Y(_1438_) );
	OR2X2 OR2X2_10 ( .A(_1437_), .B(_1438_), .Y(_1439_) );
	AOI21X1 AOI21X1_26 ( .A(dst_reg_1_), .B(_1436_), .C(_1439_), .Y(_1440_) );
	OAI22X1 OAI22X1_11 ( .A(_962__bF_buf3), .B(_1270_), .C(_957__bF_buf4), .D(_1076_), .Y(_1441_) );
	AOI21X1 AOI21X1_27 ( .A(_1119_), .B(_1270_), .C(_957__bF_buf3), .Y(_1442_) );
	NOR2X1 NOR2X1_112 ( .A(_1441_), .B(_1442_), .Y(_1443_) );
	OAI22X1 OAI22X1_12 ( .A(_1027_), .B(_962__bF_buf2), .C(_937__bF_buf1), .D(_1051_), .Y(_1444_) );
	AOI21X1 AOI21X1_28 ( .A(_963_), .B(_1046_), .C(_1444_), .Y(_1445_) );
	NAND3X1 NAND3X1_63 ( .A(_1408_), .B(_1080_), .C(_1012_), .Y(_1446_) );
	INVX1 INVX1_53 ( .A(_1446_), .Y(_1447_) );
	NAND3X1 NAND3X1_64 ( .A(_1445_), .B(_1443_), .C(_1447_), .Y(_1448_) );
	OAI21X1 OAI21X1_116 ( .A(_937__bF_buf0), .B(_1270_), .C(src_reg_1_), .Y(_1449_) );
	OAI21X1 OAI21X1_117 ( .A(_1449_), .B(_1448_), .C(_1440_), .Y(_1450_) );
	INVX1 INVX1_54 ( .A(AXYS_0__0_), .Y(_1451_) );
	AOI22X1 AOI22X1_13 ( .A(_1124_), .B(_882__bF_buf5), .C(_956_), .D(_1046_), .Y(_1452_) );
	NOR3X1 NOR3X1_13 ( .A(state_0_), .B(_1054_), .C(_948_), .Y(_1453_) );
	AOI22X1 AOI22X1_14 ( .A(_956_), .B(_1453_), .C(_947_), .D(_1046_), .Y(_1454_) );
	NAND3X1 NAND3X1_65 ( .A(_1012_), .B(_1454_), .C(_1452_), .Y(_1455_) );
	AOI22X1 AOI22X1_15 ( .A(_950_), .B(_956_), .C(_882__bF_buf4), .D(_1043_), .Y(_1456_) );
	OAI21X1 OAI21X1_118 ( .A(_972_), .B(_1124_), .C(_947_), .Y(_1457_) );
	NAND3X1 NAND3X1_66 ( .A(_1456_), .B(_1406_), .C(_1457_), .Y(_1458_) );
	NOR2X1 NOR2X1_113 ( .A(_1458_), .B(_1455_), .Y(_1459_) );
	OAI21X1 OAI21X1_119 ( .A(_937__bF_buf4), .B(_1270_), .C(src_reg_0_), .Y(_1460_) );
	NOR3X1 NOR3X1_14 ( .A(_1460_), .B(_1438_), .C(_1437_), .Y(_1461_) );
	INVX1 INVX1_55 ( .A(_1461_), .Y(_1462_) );
	NAND2X1 NAND2X1_99 ( .A(dst_reg_0_), .B(_1436_), .Y(_1463_) );
	OAI21X1 OAI21X1_120 ( .A(_1438_), .B(_1437_), .C(index_y), .Y(_1464_) );
	AND2X2 AND2X2_25 ( .A(_1464_), .B(_1463_), .Y(_1465_) );
	NAND3X1 NAND3X1_67 ( .A(_1462_), .B(_1465_), .C(_1459_), .Y(_1466_) );
	NAND2X1 NAND2X1_100 ( .A(AXYS_1__0_), .B(_1466__bF_buf4), .Y(_1467_) );
	OAI21X1 OAI21X1_121 ( .A(_1451_), .B(_1466__bF_buf3), .C(_1467_), .Y(_1468_) );
	NAND2X1 NAND2X1_101 ( .A(_1463_), .B(_1464_), .Y(_1469_) );
	NOR3X1 NOR3X1_15 ( .A(_1461_), .B(_1469_), .C(_1448_), .Y(_1470_) );
	NOR2X1 NOR2X1_114 ( .A(AXYS_3__0_), .B(_1470_), .Y(_1471_) );
	NOR2X1 NOR2X1_115 ( .A(AXYS_2__0_), .B(_1466__bF_buf2), .Y(_1472_) );
	OAI21X1 OAI21X1_122 ( .A(_1472_), .B(_1471_), .C(_1450_), .Y(_1473_) );
	OAI21X1 OAI21X1_123 ( .A(_1450_), .B(_1468_), .C(_1473_), .Y(_1474_) );
	OAI21X1 OAI21X1_124 ( .A(_957__bF_buf2), .B(_936__bF_buf3), .C(_1080_), .Y(_1475_) );
	OR2X2 OR2X2_11 ( .A(_1409_), .B(_1475_), .Y(_1476_) );
	NOR2X1 NOR2X1_116 ( .A(_1437_), .B(_1476_), .Y(_1477_) );
	INVX1 INVX1_56 ( .A(_1477_), .Y(_1478_) );
	INVX4 INVX4_9 ( .A(_1062_), .Y(_1479_) );
	INVX2 INVX2_21 ( .A(_1198_), .Y(_1480_) );
	NAND3X1 NAND3X1_68 ( .A(_1107_), .B(_1480_), .C(_1479_), .Y(_1481_) );
	NOR2X1 NOR2X1_117 ( .A(_1481_), .B(_1380_), .Y(_1482_) );
	NOR2X1 NOR2X1_118 ( .A(_1274_), .B(_1085_), .Y(_1483_) );
	NAND3X1 NAND3X1_69 ( .A(_1398_), .B(_1483_), .C(_1482_), .Y(_1484_) );
	NOR2X1 NOR2X1_119 ( .A(_1478_), .B(_1484_), .Y(_1485_) );
	OAI21X1 OAI21X1_125 ( .A(_1485_), .B(_1474_), .C(_1435_), .Y(AI_0_) );
	NAND3X1 NAND3X1_70 ( .A(ABH_1_), .B(_882__bF_buf3), .C(_1034__bF_buf2), .Y(_1486_) );
	OAI21X1 OAI21X1_126 ( .A(_1419_), .B(_1432_), .C(_1486_), .Y(_1487_) );
	AOI21X1 AOI21X1_29 ( .A(_1430_), .B(ADD_1_), .C(_1487_), .Y(_1488_) );
	INVX8 INVX8_5 ( .A(_1450_), .Y(_1489_) );
	INVX1 INVX1_57 ( .A(AXYS_0__1_), .Y(_1490_) );
	NOR2X1 NOR2X1_120 ( .A(_1490_), .B(_1466__bF_buf1), .Y(_1491_) );
	INVX1 INVX1_58 ( .A(AXYS_2__1_), .Y(_1492_) );
	NAND2X1 NAND2X1_102 ( .A(AXYS_3__1_), .B(_1466__bF_buf0), .Y(_1493_) );
	OAI21X1 OAI21X1_127 ( .A(_1492_), .B(_1466__bF_buf4), .C(_1493_), .Y(_1494_) );
	INVX1 INVX1_59 ( .A(AXYS_1__1_), .Y(_1495_) );
	OAI21X1 OAI21X1_128 ( .A(_1495_), .B(_1470_), .C(_1489_), .Y(_1496_) );
	OAI22X1 OAI22X1_13 ( .A(_1491_), .B(_1496_), .C(_1489_), .D(_1494_), .Y(_1497_) );
	OAI21X1 OAI21X1_129 ( .A(_1485_), .B(_1497_), .C(_1488_), .Y(AI_1_) );
	NAND3X1 NAND3X1_71 ( .A(ABH_2_), .B(_882__bF_buf2), .C(_1034__bF_buf1), .Y(_1498_) );
	OAI21X1 OAI21X1_130 ( .A(_905_), .B(_1432_), .C(_1498_), .Y(_1499_) );
	AOI21X1 AOI21X1_30 ( .A(_1430_), .B(ADD_2_), .C(_1499_), .Y(_1500_) );
	INVX1 INVX1_60 ( .A(AXYS_0__2_), .Y(_1501_) );
	NAND2X1 NAND2X1_103 ( .A(AXYS_1__2_), .B(_1466__bF_buf3), .Y(_1502_) );
	OAI21X1 OAI21X1_131 ( .A(_1501_), .B(_1466__bF_buf2), .C(_1502_), .Y(_1503_) );
	NOR2X1 NOR2X1_121 ( .A(AXYS_3__2_), .B(_1470_), .Y(_1504_) );
	NOR2X1 NOR2X1_122 ( .A(AXYS_2__2_), .B(_1466__bF_buf1), .Y(_1505_) );
	OAI21X1 OAI21X1_132 ( .A(_1505_), .B(_1504_), .C(_1450_), .Y(_1506_) );
	OAI21X1 OAI21X1_133 ( .A(_1450_), .B(_1503_), .C(_1506_), .Y(_1507_) );
	OAI21X1 OAI21X1_134 ( .A(_1485_), .B(_1507_), .C(_1500_), .Y(AI_2_) );
	NAND3X1 NAND3X1_72 ( .A(ABH_3_), .B(_882__bF_buf1), .C(_1034__bF_buf0), .Y(_1508_) );
	OAI21X1 OAI21X1_135 ( .A(_1095_), .B(_1432_), .C(_1508_), .Y(_1509_) );
	AOI21X1 AOI21X1_31 ( .A(_1430_), .B(ADD_3_), .C(_1509_), .Y(_1511_) );
	INVX1 INVX1_61 ( .A(AXYS_0__3_), .Y(_1512_) );
	NOR2X1 NOR2X1_123 ( .A(_1512_), .B(_1466__bF_buf0), .Y(_1514_) );
	INVX1 INVX1_62 ( .A(AXYS_2__3_), .Y(_1515_) );
	NAND2X1 NAND2X1_104 ( .A(AXYS_3__3_), .B(_1466__bF_buf4), .Y(_1517_) );
	OAI21X1 OAI21X1_136 ( .A(_1515_), .B(_1466__bF_buf3), .C(_1517_), .Y(_1518_) );
	INVX1 INVX1_63 ( .A(AXYS_1__3_), .Y(_1520_) );
	OAI21X1 OAI21X1_137 ( .A(_1520_), .B(_1470_), .C(_1489_), .Y(_1521_) );
	OAI22X1 OAI22X1_14 ( .A(_1514_), .B(_1521_), .C(_1489_), .D(_1518_), .Y(_1523_) );
	OAI21X1 OAI21X1_138 ( .A(_1485_), .B(_1523_), .C(_1511_), .Y(AI_3_) );
	INVX2 INVX2_22 ( .A(ABH_4_), .Y(_1525_) );
	OAI22X1 OAI22X1_15 ( .A(_1525_), .B(_1064_), .C(_891_), .D(_1432_), .Y(_1526_) );
	AOI21X1 AOI21X1_32 ( .A(_1430_), .B(ADD_4_), .C(_1526_), .Y(_1528_) );
	INVX1 INVX1_64 ( .A(AXYS_0__4_), .Y(_1529_) );
	NAND2X1 NAND2X1_105 ( .A(AXYS_1__4_), .B(_1466__bF_buf2), .Y(_1531_) );
	OAI21X1 OAI21X1_139 ( .A(_1529_), .B(_1466__bF_buf1), .C(_1531_), .Y(_1532_) );
	NOR2X1 NOR2X1_124 ( .A(AXYS_3__4_), .B(_1470_), .Y(_1533_) );
	NOR2X1 NOR2X1_125 ( .A(AXYS_2__4_), .B(_1466__bF_buf0), .Y(_1534_) );
	OAI21X1 OAI21X1_140 ( .A(_1534_), .B(_1533_), .C(_1450_), .Y(_1535_) );
	OAI21X1 OAI21X1_141 ( .A(_1450_), .B(_1532_), .C(_1535_), .Y(_41_) );
	OAI21X1 OAI21X1_142 ( .A(_1485_), .B(_41_), .C(_1528_), .Y(AI_4_) );
	INVX1 INVX1_65 ( .A(ABH_5_), .Y(_42_) );
	OAI22X1 OAI22X1_16 ( .A(_42_), .B(_1064_), .C(_1424_), .D(_1432_), .Y(_43_) );
	AOI21X1 AOI21X1_33 ( .A(_1430_), .B(ADD_5_), .C(_43_), .Y(_44_) );
	INVX1 INVX1_66 ( .A(AXYS_0__5_), .Y(_45_) );
	NAND2X1 NAND2X1_106 ( .A(AXYS_1__5_), .B(_1466__bF_buf4), .Y(_46_) );
	OAI21X1 OAI21X1_143 ( .A(_45_), .B(_1466__bF_buf3), .C(_46_), .Y(_47_) );
	NOR2X1 NOR2X1_126 ( .A(AXYS_3__5_), .B(_1470_), .Y(_48_) );
	NOR2X1 NOR2X1_127 ( .A(AXYS_2__5_), .B(_1466__bF_buf2), .Y(_49_) );
	OAI21X1 OAI21X1_144 ( .A(_49_), .B(_48_), .C(_1450_), .Y(_50_) );
	OAI21X1 OAI21X1_145 ( .A(_1450_), .B(_47_), .C(_50_), .Y(_51_) );
	OAI21X1 OAI21X1_146 ( .A(_1485_), .B(_51_), .C(_44_), .Y(AI_5_) );
	INVX2 INVX2_23 ( .A(ABH_6_), .Y(_52_) );
	OAI22X1 OAI22X1_17 ( .A(_52_), .B(_1064_), .C(_1260_), .D(_1432_), .Y(_53_) );
	AOI21X1 AOI21X1_34 ( .A(_1430_), .B(ADD_6_), .C(_53_), .Y(_54_) );
	INVX1 INVX1_67 ( .A(AXYS_0__6_), .Y(_55_) );
	NAND2X1 NAND2X1_107 ( .A(AXYS_1__6_), .B(_1466__bF_buf1), .Y(_56_) );
	OAI21X1 OAI21X1_147 ( .A(_55_), .B(_1466__bF_buf0), .C(_56_), .Y(_57_) );
	NOR2X1 NOR2X1_128 ( .A(AXYS_3__6_), .B(_1470_), .Y(_58_) );
	NOR2X1 NOR2X1_129 ( .A(AXYS_2__6_), .B(_1466__bF_buf4), .Y(_59_) );
	OAI21X1 OAI21X1_148 ( .A(_59_), .B(_58_), .C(_1450_), .Y(_60_) );
	OAI21X1 OAI21X1_149 ( .A(_1450_), .B(_57_), .C(_60_), .Y(_61_) );
	OAI21X1 OAI21X1_150 ( .A(_1485_), .B(_61_), .C(_54_), .Y(AI_6_) );
	INVX2 INVX2_24 ( .A(ABH_7_), .Y(_62_) );
	OAI22X1 OAI22X1_18 ( .A(_62_), .B(_1064_), .C(_925_), .D(_1432_), .Y(_63_) );
	AOI21X1 AOI21X1_35 ( .A(_1430_), .B(ADD_7_), .C(_63_), .Y(_64_) );
	INVX1 INVX1_68 ( .A(AXYS_0__7_), .Y(_65_) );
	NOR2X1 NOR2X1_130 ( .A(_65_), .B(_1466__bF_buf3), .Y(_66_) );
	INVX1 INVX1_69 ( .A(AXYS_2__7_), .Y(_67_) );
	NAND2X1 NAND2X1_108 ( .A(AXYS_3__7_), .B(_1466__bF_buf2), .Y(_69_) );
	OAI21X1 OAI21X1_151 ( .A(_67_), .B(_1466__bF_buf1), .C(_69_), .Y(_70_) );
	INVX1 INVX1_70 ( .A(AXYS_1__7_), .Y(_72_) );
	OAI21X1 OAI21X1_152 ( .A(_72_), .B(_1470_), .C(_1489_), .Y(_73_) );
	OAI22X1 OAI22X1_19 ( .A(_66_), .B(_73_), .C(_1489_), .D(_70_), .Y(_75_) );
	OAI21X1 OAI21X1_153 ( .A(_1485_), .B(_75_), .C(_64_), .Y(AI_7_) );
	INVX1 INVX1_71 ( .A(op_0_), .Y(_77_) );
	INVX2 INVX2_25 ( .A(_1379_), .Y(_78_) );
	OAI21X1 OAI21X1_154 ( .A(_972_), .B(_954_), .C(_882__bF_buf0), .Y(_80_) );
	NAND2X1 NAND2X1_109 ( .A(_80_), .B(_78_), .Y(_81_) );
	OAI21X1 OAI21X1_155 ( .A(_77_), .B(_78_), .C(_81_), .Y(ALU_op_0_) );
	INVX1 INVX1_72 ( .A(op_1_), .Y(_83_) );
	OAI21X1 OAI21X1_156 ( .A(_83_), .B(_78_), .C(_81_), .Y(ALU_op_1_) );
	INVX1 INVX1_73 ( .A(backwards), .Y(_85_) );
	OAI21X1 OAI21X1_157 ( .A(_957__bF_buf1), .B(_1076_), .C(_1452_), .Y(_87_) );
	OAI21X1 OAI21X1_158 ( .A(_962__bF_buf1), .B(_1051_), .C(_1193_), .Y(_88_) );
	INVX4 INVX4_10 ( .A(_88_), .Y(_89_) );
	OAI21X1 OAI21X1_159 ( .A(_937__bF_buf3), .B(_1061_), .C(_89_), .Y(_90_) );
	NOR2X1 NOR2X1_131 ( .A(_87_), .B(_90_), .Y(_91_) );
	INVX1 INVX1_74 ( .A(_91_), .Y(_92_) );
	AOI21X1 AOI21X1_36 ( .A(op_2_), .B(_1379_), .C(_92_), .Y(_93_) );
	OAI21X1 OAI21X1_160 ( .A(_85_), .B(_1064_), .C(_93_), .Y(ALU_op_2_) );
	INVX1 INVX1_75 ( .A(op_3_), .Y(_94_) );
	NOR2X1 NOR2X1_132 ( .A(_94_), .B(_78_), .Y(ALU_op_3_) );
	INVX2 INVX2_26 ( .A(_959_), .Y(_95_) );
	NOR2X1 NOR2X1_133 ( .A(_1020_), .B(_967_), .Y(_96_) );
	OAI21X1 OAI21X1_161 ( .A(_955_), .B(_936__bF_buf2), .C(_96_), .Y(_97_) );
	OAI21X1 OAI21X1_162 ( .A(_943_), .B(_97_), .C(store), .Y(_98_) );
	NAND3X1 NAND3X1_73 ( .A(_95_), .B(_98_), .C(_91_), .Y(_1538_) );
	OAI21X1 OAI21X1_163 ( .A(_957__bF_buf0), .B(_958_), .C(_91_), .Y(_99_) );
	AND2X2 AND2X2_26 ( .A(_1198_), .B(php), .Y(_100_) );
	OAI21X1 OAI21X1_164 ( .A(_1194_), .B(_100_), .C(C), .Y(_101_) );
	INVX1 INVX1_76 ( .A(PC_8_), .Y(_102_) );
	OAI22X1 OAI22X1_20 ( .A(_102_), .B(_1452_), .C(_1402_), .D(_89_), .Y(_103_) );
	OAI21X1 OAI21X1_165 ( .A(php), .B(_1480_), .C(_95_), .Y(_104_) );
	AOI21X1 AOI21X1_37 ( .A(ADD_0_), .B(_104_), .C(_103_), .Y(_105_) );
	AND2X2 AND2X2_27 ( .A(_105_), .B(_101_), .Y(_106_) );
	OAI21X1 OAI21X1_166 ( .A(_99_), .B(_1474_), .C(_106_), .Y(_1537__0_) );
	INVX2 INVX2_27 ( .A(PC_9_), .Y(_107_) );
	NOR2X1 NOR2X1_134 ( .A(_99_), .B(_1497_), .Y(_108_) );
	MUX2X1 MUX2X1_8 ( .A(Z), .B(ADD_1_), .S(php), .Y(_109_) );
	OAI22X1 OAI22X1_21 ( .A(_1174_), .B(_1057__bF_buf0), .C(_109_), .D(_1480_), .Y(_110_) );
	AOI21X1 AOI21X1_38 ( .A(ADD_1_), .B(_959_), .C(_110_), .Y(_111_) );
	OAI21X1 OAI21X1_167 ( .A(_1418_), .B(_89_), .C(_111_), .Y(_112_) );
	NOR2X1 NOR2X1_135 ( .A(_112_), .B(_108_), .Y(_113_) );
	OAI21X1 OAI21X1_168 ( .A(_107_), .B(_1452_), .C(_113_), .Y(_1537__1_) );
	INVX2 INVX2_28 ( .A(PC_10_), .Y(_114_) );
	INVX4 INVX4_11 ( .A(ADD_2_), .Y(_115_) );
	NAND2X1 NAND2X1_110 ( .A(php), .B(I), .Y(_116_) );
	OAI21X1 OAI21X1_169 ( .A(php), .B(_115_), .C(_116_), .Y(_117_) );
	OAI22X1 OAI22X1_22 ( .A(_892_), .B(_1057__bF_buf3), .C(_115_), .D(_95_), .Y(_118_) );
	AOI21X1 AOI21X1_39 ( .A(_1198_), .B(_117_), .C(_118_), .Y(_119_) );
	OAI21X1 OAI21X1_170 ( .A(_114_), .B(_1452_), .C(_119_), .Y(_120_) );
	AOI21X1 AOI21X1_40 ( .A(PC_2_), .B(_88_), .C(_120_), .Y(_121_) );
	OAI21X1 OAI21X1_171 ( .A(_99_), .B(_1507_), .C(_121_), .Y(_1537__2_) );
	INVX2 INVX2_29 ( .A(PC_11_), .Y(_122_) );
	NOR2X1 NOR2X1_136 ( .A(_99_), .B(_1523_), .Y(_123_) );
	INVX1 INVX1_77 ( .A(D), .Y(_124_) );
	MUX2X1 MUX2X1_9 ( .A(D), .B(ADD_3_), .S(php), .Y(_125_) );
	OAI22X1 OAI22X1_23 ( .A(_124_), .B(_1057__bF_buf2), .C(_125_), .D(_1480_), .Y(_126_) );
	AOI21X1 AOI21X1_41 ( .A(ADD_3_), .B(_959_), .C(_126_), .Y(_127_) );
	OAI21X1 OAI21X1_172 ( .A(_1421_), .B(_89_), .C(_127_), .Y(_128_) );
	NOR2X1 NOR2X1_137 ( .A(_128_), .B(_123_), .Y(_129_) );
	OAI21X1 OAI21X1_173 ( .A(_122_), .B(_1452_), .C(_129_), .Y(_1537__3_) );
	OAI22X1 OAI22X1_24 ( .A(_959_), .B(_1198_), .C(ADD_4_), .D(_100_), .Y(_130_) );
	INVX2 INVX2_30 ( .A(PC_12_), .Y(_131_) );
	OAI22X1 OAI22X1_25 ( .A(_895_), .B(_1057__bF_buf1), .C(_131_), .D(_1452_), .Y(_132_) );
	AOI21X1 AOI21X1_42 ( .A(PC_4_), .B(_88_), .C(_132_), .Y(_133_) );
	AND2X2 AND2X2_28 ( .A(_133_), .B(_130_), .Y(_134_) );
	OAI21X1 OAI21X1_174 ( .A(_99_), .B(_41_), .C(_134_), .Y(_1537__4_) );
	INVX1 INVX1_78 ( .A(PC_13_), .Y(_135_) );
	NOR2X1 NOR2X1_138 ( .A(_1194_), .B(_100_), .Y(_136_) );
	OAI21X1 OAI21X1_175 ( .A(_135_), .B(_1452_), .C(_136_), .Y(_137_) );
	OAI21X1 OAI21X1_176 ( .A(_1198_), .B(_959_), .C(ADD_5_), .Y(_138_) );
	OAI21X1 OAI21X1_177 ( .A(_1423_), .B(_89_), .C(_138_), .Y(_139_) );
	NOR2X1 NOR2X1_139 ( .A(_137_), .B(_139_), .Y(_140_) );
	OAI21X1 OAI21X1_178 ( .A(_99_), .B(_51_), .C(_140_), .Y(_1537__5_) );
	OAI21X1 OAI21X1_179 ( .A(_1194_), .B(_100_), .C(V), .Y(_141_) );
	INVX1 INVX1_79 ( .A(PC_14_), .Y(_142_) );
	OAI22X1 OAI22X1_26 ( .A(_142_), .B(_1452_), .C(_1425_), .D(_89_), .Y(_143_) );
	AOI21X1 AOI21X1_43 ( .A(ADD_6_), .B(_104_), .C(_143_), .Y(_144_) );
	AND2X2 AND2X2_29 ( .A(_144_), .B(_141_), .Y(_145_) );
	OAI21X1 OAI21X1_180 ( .A(_99_), .B(_61_), .C(_145_), .Y(_1537__6_) );
	OAI21X1 OAI21X1_181 ( .A(_1194_), .B(_100_), .C(N), .Y(_146_) );
	INVX1 INVX1_80 ( .A(PC_15_), .Y(_147_) );
	OAI22X1 OAI22X1_27 ( .A(_147_), .B(_1452_), .C(_1426_), .D(_89_), .Y(_148_) );
	AOI21X1 AOI21X1_44 ( .A(ADD_7_), .B(_104_), .C(_148_), .Y(_149_) );
	AND2X2 AND2X2_30 ( .A(_149_), .B(_146_), .Y(_150_) );
	OAI21X1 OAI21X1_182 ( .A(_99_), .B(_75_), .C(_150_), .Y(_1537__7_) );
	INVX2 INVX2_31 ( .A(adc_sbc), .Y(_151_) );
	NOR2X1 NOR2X1_140 ( .A(_124_), .B(_151_), .Y(_14_) );
	INVX1 INVX1_81 ( .A(adc_bcd), .Y(_152_) );
	NOR2X1 NOR2X1_141 ( .A(_152_), .B(_978_), .Y(ALU_BCD) );
	INVX4 INVX4_12 ( .A(reset), .Y(_1214_) );
	INVX1 INVX1_82 ( .A(res), .Y(_155_) );
	OAI21X1 OAI21X1_183 ( .A(_155_), .B(_1436_), .C(_1214_), .Y(_31_) );
	NAND2X1 NAND2X1_111 ( .A(plp), .B(_1436_), .Y(_157_) );
	INVX2 INVX2_32 ( .A(plp), .Y(_158_) );
	OAI21X1 OAI21X1_184 ( .A(_158_), .B(_885__bF_buf1), .C(I), .Y(_160_) );
	OAI21X1 OAI21X1_185 ( .A(_115_), .B(_157_), .C(_160_), .Y(_161_) );
	NOR2X1 NOR2X1_142 ( .A(_1219_), .B(_161_), .Y(_163_) );
	INVX1 INVX1_83 ( .A(_1219_), .Y(_164_) );
	INVX1 INVX1_84 ( .A(sei), .Y(_166_) );
	AOI21X1 AOI21X1_45 ( .A(_892_), .B(_166_), .C(cli), .Y(_167_) );
	OAI21X1 OAI21X1_186 ( .A(_167_), .B(_164_), .C(_1392_), .Y(_169_) );
	AOI21X1 AOI21X1_46 ( .A(_1038_), .B(DIMUX_2_), .C(_1052_), .Y(_170_) );
	OAI21X1 OAI21X1_187 ( .A(_169_), .B(_163_), .C(_170_), .Y(_6_) );
	AND2X2 AND2X2_31 ( .A(_1379_), .B(shift_right), .Y(ALU_right) );
	NAND2X1 NAND2X1_112 ( .A(load_reg), .B(_158_), .Y(_172_) );
	OAI21X1 OAI21X1_188 ( .A(_885__bF_buf0), .B(_172_), .C(_1456_), .Y(_173_) );
	OAI21X1 OAI21X1_189 ( .A(_972_), .B(_1046_), .C(_956_), .Y(_174_) );
	NAND2X1 NAND2X1_113 ( .A(_1457_), .B(_174_), .Y(_175_) );
	OAI21X1 OAI21X1_190 ( .A(_173_), .B(_175_), .C(RDY_bF_buf6), .Y(_176_) );
	INVX1 INVX1_85 ( .A(_176_), .Y(_177_) );
	NAND2X1 NAND2X1_114 ( .A(_177_), .B(_1470_), .Y(_178_) );
	NOR2X1 NOR2X1_143 ( .A(_1450_), .B(_178_), .Y(_179_) );
	OAI21X1 OAI21X1_191 ( .A(_962__bF_buf0), .B(_1061_), .C(ADD_0_), .Y(_180_) );
	OAI21X1 OAI21X1_192 ( .A(_1403_), .B(_1479_), .C(_180_), .Y(_181_) );
	NAND2X1 NAND2X1_115 ( .A(_181_), .B(_179_), .Y(_182_) );
	OAI21X1 OAI21X1_193 ( .A(_1451_), .B(_179_), .C(_182_), .Y(_1328_) );
	NAND3X1 NAND3X1_74 ( .A(adc_bcd), .B(adj_bcd), .C(ALU_HC), .Y(_183_) );
	NAND2X1 NAND2X1_116 ( .A(adj_bcd), .B(_152_), .Y(_184_) );
	OAI21X1 OAI21X1_194 ( .A(ALU_HC), .B(_184_), .C(_183_), .Y(_185_) );
	NAND2X1 NAND2X1_117 ( .A(ADD_1_), .B(_185_), .Y(_186_) );
	INVX1 INVX1_86 ( .A(_186_), .Y(_187_) );
	NOR2X1 NOR2X1_144 ( .A(_1062_), .B(_187_), .Y(_188_) );
	OAI21X1 OAI21X1_195 ( .A(ADD_1_), .B(_185_), .C(_188_), .Y(_189_) );
	OAI21X1 OAI21X1_196 ( .A(_1419_), .B(_1479_), .C(_189_), .Y(_190_) );
	NAND2X1 NAND2X1_118 ( .A(_190_), .B(_179_), .Y(_191_) );
	OAI21X1 OAI21X1_197 ( .A(_1490_), .B(_179_), .C(_191_), .Y(_1345_) );
	XNOR2X1 XNOR2X1_2 ( .A(_183_), .B(ADD_2_), .Y(_192_) );
	NOR2X1 NOR2X1_145 ( .A(_192_), .B(_187_), .Y(_193_) );
	NAND2X1 NAND2X1_119 ( .A(_192_), .B(_187_), .Y(_194_) );
	OAI21X1 OAI21X1_198 ( .A(_962__bF_buf4), .B(_1061_), .C(_194_), .Y(_195_) );
	OAI22X1 OAI22X1_28 ( .A(_905_), .B(_1479_), .C(_193_), .D(_195_), .Y(_196_) );
	NAND2X1 NAND2X1_120 ( .A(_196_), .B(_179_), .Y(_197_) );
	OAI21X1 OAI21X1_199 ( .A(_1501_), .B(_179_), .C(_197_), .Y(_1352_) );
	OAI21X1 OAI21X1_200 ( .A(_115_), .B(_183_), .C(_194_), .Y(_198_) );
	INVX2 INVX2_33 ( .A(ADD_3_), .Y(_199_) );
	NOR2X1 NOR2X1_146 ( .A(ALU_HC), .B(_184_), .Y(_200_) );
	XNOR2X1 XNOR2X1_3 ( .A(_200_), .B(_199_), .Y(_201_) );
	XNOR2X1 XNOR2X1_4 ( .A(_198_), .B(_201_), .Y(_202_) );
	NAND2X1 NAND2X1_121 ( .A(DIMUX_3_), .B(_1062_), .Y(_203_) );
	OAI21X1 OAI21X1_201 ( .A(_1062_), .B(_202_), .C(_203_), .Y(_204_) );
	NAND2X1 NAND2X1_122 ( .A(_179_), .B(_204_), .Y(_205_) );
	OAI21X1 OAI21X1_202 ( .A(_1512_), .B(_179_), .C(_205_), .Y(_1359_) );
	OAI21X1 OAI21X1_203 ( .A(_962__bF_buf3), .B(_1061_), .C(ADD_4_), .Y(_206_) );
	OAI21X1 OAI21X1_204 ( .A(_891_), .B(_1479_), .C(_206_), .Y(_207_) );
	NAND2X1 NAND2X1_123 ( .A(_207_), .B(_179_), .Y(_208_) );
	OAI21X1 OAI21X1_205 ( .A(_1529_), .B(_179_), .C(_208_), .Y(_1363_) );
	INVX2 INVX2_34 ( .A(ADD_5_), .Y(_209_) );
	NAND3X1 NAND3X1_75 ( .A(ALU_CO), .B(adc_bcd), .C(adj_bcd), .Y(_210_) );
	INVX1 INVX1_87 ( .A(_210_), .Y(_211_) );
	NOR2X1 NOR2X1_147 ( .A(ALU_CO), .B(_184_), .Y(_212_) );
	NOR2X1 NOR2X1_148 ( .A(_211_), .B(_212_), .Y(_213_) );
	NAND2X1 NAND2X1_124 ( .A(_209_), .B(_213_), .Y(_214_) );
	NOR2X1 NOR2X1_149 ( .A(_209_), .B(_213_), .Y(_215_) );
	NOR2X1 NOR2X1_150 ( .A(_1062_), .B(_215_), .Y(_216_) );
	AOI22X1 AOI22X1_16 ( .A(DIMUX_5_), .B(_1062_), .C(_214_), .D(_216_), .Y(_217_) );
	MUX2X1 MUX2X1_10 ( .A(_217_), .B(_45_), .S(_179_), .Y(_1375_) );
	XNOR2X1 XNOR2X1_5 ( .A(_210_), .B(ADD_6_), .Y(_218_) );
	NAND2X1 NAND2X1_125 ( .A(_218_), .B(_215_), .Y(_219_) );
	OR2X2 OR2X2_12 ( .A(_215_), .B(_218_), .Y(_220_) );
	NAND3X1 NAND3X1_76 ( .A(_1479_), .B(_219_), .C(_220_), .Y(_221_) );
	OAI21X1 OAI21X1_206 ( .A(_1260_), .B(_1479_), .C(_221_), .Y(_222_) );
	NAND2X1 NAND2X1_126 ( .A(_222_), .B(_179_), .Y(_223_) );
	OAI21X1 OAI21X1_207 ( .A(_55_), .B(_179_), .C(_223_), .Y(_1381_) );
	INVX2 INVX2_35 ( .A(ADD_6_), .Y(_224_) );
	OAI21X1 OAI21X1_208 ( .A(_224_), .B(_210_), .C(_219_), .Y(_225_) );
	XNOR2X1 XNOR2X1_6 ( .A(_212_), .B(ADD_7_), .Y(_226_) );
	XNOR2X1 XNOR2X1_7 ( .A(_225_), .B(_226_), .Y(_227_) );
	OAI21X1 OAI21X1_209 ( .A(_962__bF_buf2), .B(_1061_), .C(_227_), .Y(_228_) );
	OAI21X1 OAI21X1_210 ( .A(_925_), .B(_1479_), .C(_228_), .Y(_229_) );
	NAND2X1 NAND2X1_127 ( .A(_179_), .B(_229_), .Y(_230_) );
	OAI21X1 OAI21X1_211 ( .A(_65_), .B(_179_), .C(_230_), .Y(_1389_) );
	INVX1 INVX1_88 ( .A(NMI_1), .Y(_231_) );
	NAND3X1 NAND3X1_77 ( .A(NMI), .B(_894_), .C(_231_), .Y(_232_) );
	OAI21X1 OAI21X1_212 ( .A(_894_), .B(_1052_), .C(_232_), .Y(_7_) );
	NAND2X1 NAND2X1_128 ( .A(cond_code_0_), .B(_881__bF_buf2), .Y(_233_) );
	OAI21X1 OAI21X1_213 ( .A(_881__bF_buf1), .B(_1162_), .C(_233_), .Y(_22__0_) );
	NAND2X1 NAND2X1_129 ( .A(cond_code_1_), .B(_881__bF_buf0), .Y(_234_) );
	OAI21X1 OAI21X1_214 ( .A(_881__bF_buf7), .B(_1008_), .C(_234_), .Y(_22__1_) );
	NAND2X1 NAND2X1_130 ( .A(cond_code_2_), .B(_881__bF_buf6), .Y(_235_) );
	OAI21X1 OAI21X1_215 ( .A(_881__bF_buf5), .B(_1092_), .C(_235_), .Y(_22__2_) );
	NAND2X1 NAND2X1_131 ( .A(_886__bF_buf4), .B(_1100_), .Y(_236_) );
	NAND2X1 NAND2X1_132 ( .A(_1008_), .B(_928_), .Y(_237_) );
	INVX1 INVX1_89 ( .A(_237_), .Y(_238_) );
	NAND2X1 NAND2X1_133 ( .A(_1003_), .B(_238_), .Y(_239_) );
	NOR2X1 NOR2X1_151 ( .A(_924_), .B(_239_), .Y(_240_) );
	INVX1 INVX1_90 ( .A(_240_), .Y(_241_) );
	OAI21X1 OAI21X1_216 ( .A(_881__bF_buf4), .B(_885__bF_buf4), .C(clv), .Y(_242_) );
	OAI21X1 OAI21X1_217 ( .A(_236_), .B(_241_), .C(_242_), .Y(_20_) );
	NAND2X1 NAND2X1_134 ( .A(_1003_), .B(_1206_), .Y(_243_) );
	NAND2X1 NAND2X1_135 ( .A(_1169_), .B(_1100_), .Y(_244_) );
	OAI22X1 OAI22X1_29 ( .A(_166_), .B(_886__bF_buf3), .C(_243_), .D(_244_), .Y(_35_) );
	OAI21X1 OAI21X1_218 ( .A(_881__bF_buf3), .B(_885__bF_buf3), .C(cli), .Y(_245_) );
	OAI21X1 OAI21X1_219 ( .A(_910__bF_buf3), .B(_1002_), .C(_1206_), .Y(_246_) );
	OAI21X1 OAI21X1_220 ( .A(_246_), .B(_244_), .C(_245_), .Y(_19_) );
	OAI21X1 OAI21X1_221 ( .A(_881__bF_buf2), .B(_885__bF_buf2), .C(sed), .Y(_247_) );
	NOR2X1 NOR2X1_152 ( .A(_1092_), .B(_1008_), .Y(_248_) );
	NAND2X1 NAND2X1_136 ( .A(_248_), .B(_1100_), .Y(_249_) );
	OAI21X1 OAI21X1_222 ( .A(_243_), .B(_249_), .C(_247_), .Y(_34_) );
	OAI21X1 OAI21X1_223 ( .A(_881__bF_buf1), .B(_885__bF_buf1), .C(cld), .Y(_250_) );
	OAI21X1 OAI21X1_224 ( .A(_246_), .B(_249_), .C(_250_), .Y(_18_) );
	INVX1 INVX1_91 ( .A(sec), .Y(_251_) );
	NAND2X1 NAND2X1_137 ( .A(_1165_), .B(_1100_), .Y(_252_) );
	OAI22X1 OAI22X1_30 ( .A(_251_), .B(_886__bF_buf2), .C(_243_), .D(_252_), .Y(_33_) );
	OAI21X1 OAI21X1_225 ( .A(_881__bF_buf0), .B(_885__bF_buf0), .C(clc), .Y(_253_) );
	OAI21X1 OAI21X1_226 ( .A(_246_), .B(_252_), .C(_253_), .Y(_17_) );
	OAI21X1 OAI21X1_227 ( .A(_881__bF_buf7), .B(_885__bF_buf4), .C(php), .Y(_254_) );
	OAI21X1 OAI21X1_228 ( .A(_1258_), .B(_236_), .C(_254_), .Y(_29_) );
	OAI22X1 OAI22X1_31 ( .A(_158_), .B(_886__bF_buf1), .C(_1166_), .D(_236_), .Y(_30_) );
	INVX2 INVX2_36 ( .A(bit_ins), .Y(_255_) );
	OAI21X1 OAI21X1_229 ( .A(_910__bF_buf2), .B(_913_), .C(_1148_), .Y(_256_) );
	NOR2X1 NOR2X1_153 ( .A(_256_), .B(_1166_), .Y(_257_) );
	NAND2X1 NAND2X1_138 ( .A(_886__bF_buf0), .B(_257_), .Y(_258_) );
	OAI21X1 OAI21X1_230 ( .A(_255_), .B(_886__bF_buf4), .C(_258_), .Y(_16_) );
	NAND2X1 NAND2X1_139 ( .A(_1003_), .B(_1262_), .Y(_259_) );
	NAND3X1 NAND3X1_78 ( .A(_1092_), .B(_259_), .C(_919_), .Y(_260_) );
	INVX1 INVX1_92 ( .A(_260_), .Y(_261_) );
	AOI21X1 AOI21X1_47 ( .A(_261_), .B(_1003_), .C(_1022__bF_buf2), .Y(_262_) );
	AOI22X1 AOI22X1_17 ( .A(_77_), .B(_1022__bF_buf1), .C(_261_), .D(_262_), .Y(_28__0_) );
	OAI21X1 OAI21X1_231 ( .A(_881__bF_buf6), .B(_885__bF_buf3), .C(_83_), .Y(_263_) );
	NAND2X1 NAND2X1_140 ( .A(_248_), .B(_995_), .Y(_264_) );
	INVX1 INVX1_93 ( .A(_264_), .Y(_265_) );
	INVX1 INVX1_94 ( .A(_248_), .Y(_266_) );
	NOR2X1 NOR2X1_154 ( .A(_898_), .B(_266_), .Y(_267_) );
	AOI22X1 AOI22X1_18 ( .A(_267_), .B(_1247_), .C(_1021_), .D(_265_), .Y(_268_) );
	NOR2X1 NOR2X1_155 ( .A(_1256_), .B(_237_), .Y(_269_) );
	OAI21X1 OAI21X1_232 ( .A(_910__bF_buf1), .B(_1002_), .C(_908_), .Y(_270_) );
	OAI21X1 OAI21X1_233 ( .A(_270_), .B(_1249_), .C(_1203_), .Y(_271_) );
	AOI22X1 AOI22X1_19 ( .A(_271_), .B(_248_), .C(_1100_), .D(_269_), .Y(_272_) );
	INVX1 INVX1_95 ( .A(_929_), .Y(_273_) );
	NAND3X1 NAND3X1_79 ( .A(_273_), .B(_1009_), .C(_1254_), .Y(_274_) );
	NAND3X1 NAND3X1_80 ( .A(_272_), .B(_274_), .C(_268_), .Y(_275_) );
	NOR2X1 NOR2X1_156 ( .A(_261_), .B(_257_), .Y(_276_) );
	OAI21X1 OAI21X1_234 ( .A(_1263_), .B(_1249_), .C(_276_), .Y(_277_) );
	NOR2X1 NOR2X1_157 ( .A(_275_), .B(_277_), .Y(_278_) );
	OAI21X1 OAI21X1_235 ( .A(_1164_), .B(_1249_), .C(_278_), .Y(_279_) );
	NOR2X1 NOR2X1_158 ( .A(_928_), .B(_1249_), .Y(_280_) );
	NOR2X1 NOR2X1_159 ( .A(_1022__bF_buf0), .B(_280_), .Y(_281_) );
	AND2X2 AND2X2_32 ( .A(_919_), .B(_1009_), .Y(_282_) );
	AOI21X1 AOI21X1_48 ( .A(_1092_), .B(_282_), .C(_275_), .Y(_283_) );
	NAND3X1 NAND3X1_81 ( .A(_281_), .B(_283_), .C(_279_), .Y(_284_) );
	AND2X2 AND2X2_33 ( .A(_284_), .B(_263_), .Y(_28__1_) );
	OAI21X1 OAI21X1_236 ( .A(_881__bF_buf5), .B(_885__bF_buf2), .C(op_2_), .Y(_285_) );
	OAI21X1 OAI21X1_237 ( .A(_1022__bF_buf3), .B(_278_), .C(_285_), .Y(_28__2_) );
	AOI22X1 AOI22X1_20 ( .A(_94_), .B(_1022__bF_buf2), .C(_281_), .D(_276_), .Y(_28__3_) );
	INVX1 INVX1_96 ( .A(_181_), .Y(_286_) );
	NOR2X1 NOR2X1_160 ( .A(_1489_), .B(_178_), .Y(_287_) );
	INVX4 INVX4_13 ( .A(_287_), .Y(_288_) );
	OAI21X1 OAI21X1_238 ( .A(_1489_), .B(_178_), .C(AXYS_2__0_), .Y(_289_) );
	OAI21X1 OAI21X1_239 ( .A(_286_), .B(_288_), .C(_289_), .Y(_1510_) );
	INVX1 INVX1_97 ( .A(_190_), .Y(_290_) );
	OAI21X1 OAI21X1_240 ( .A(_1489_), .B(_178_), .C(AXYS_2__1_), .Y(_291_) );
	OAI21X1 OAI21X1_241 ( .A(_290_), .B(_288_), .C(_291_), .Y(_1513_) );
	INVX1 INVX1_98 ( .A(_196_), .Y(_292_) );
	OAI21X1 OAI21X1_242 ( .A(_1489_), .B(_178_), .C(AXYS_2__2_), .Y(_293_) );
	OAI21X1 OAI21X1_243 ( .A(_292_), .B(_288_), .C(_293_), .Y(_1516_) );
	INVX1 INVX1_99 ( .A(_204_), .Y(_294_) );
	OAI21X1 OAI21X1_244 ( .A(_1489_), .B(_178_), .C(AXYS_2__3_), .Y(_295_) );
	OAI21X1 OAI21X1_245 ( .A(_288_), .B(_294_), .C(_295_), .Y(_1519_) );
	INVX1 INVX1_100 ( .A(_207_), .Y(_296_) );
	OAI21X1 OAI21X1_246 ( .A(_1489_), .B(_178_), .C(AXYS_2__4_), .Y(_297_) );
	OAI21X1 OAI21X1_247 ( .A(_296_), .B(_288_), .C(_297_), .Y(_1522_) );
	OAI21X1 OAI21X1_248 ( .A(_1489_), .B(_178_), .C(AXYS_2__5_), .Y(_298_) );
	OAI21X1 OAI21X1_249 ( .A(_217_), .B(_288_), .C(_298_), .Y(_1524_) );
	INVX1 INVX1_101 ( .A(_222_), .Y(_299_) );
	OAI21X1 OAI21X1_250 ( .A(_1489_), .B(_178_), .C(AXYS_2__6_), .Y(_300_) );
	OAI21X1 OAI21X1_251 ( .A(_299_), .B(_288_), .C(_300_), .Y(_1527_) );
	INVX1 INVX1_102 ( .A(_229_), .Y(_301_) );
	OAI21X1 OAI21X1_252 ( .A(_1489_), .B(_178_), .C(AXYS_2__7_), .Y(_302_) );
	OAI21X1 OAI21X1_253 ( .A(_288_), .B(_301_), .C(_302_), .Y(_1530_) );
	NOR2X1 NOR2X1_161 ( .A(_928_), .B(_1162_), .Y(_303_) );
	NAND2X1 NAND2X1_141 ( .A(_908_), .B(_1003_), .Y(_304_) );
	NOR2X1 NOR2X1_162 ( .A(_304_), .B(_1249_), .Y(_305_) );
	AOI22X1 AOI22X1_21 ( .A(_305_), .B(_1092_), .C(_303_), .D(_1254_), .Y(_306_) );
	OAI21X1 OAI21X1_254 ( .A(_881__bF_buf4), .B(_885__bF_buf1), .C(rotate), .Y(_307_) );
	OAI21X1 OAI21X1_255 ( .A(_1022__bF_buf1), .B(_306_), .C(_307_), .Y(_32_) );
	NOR2X1 NOR2X1_163 ( .A(_1249_), .B(_1263_), .Y(_308_) );
	INVX1 INVX1_103 ( .A(_308_), .Y(_309_) );
	OAI21X1 OAI21X1_256 ( .A(_881__bF_buf3), .B(_885__bF_buf0), .C(shift_right), .Y(_310_) );
	OAI21X1 OAI21X1_257 ( .A(_1022__bF_buf0), .B(_309_), .C(_310_), .Y(_37_) );
	AOI21X1 AOI21X1_49 ( .A(_282_), .B(_928_), .C(_1022__bF_buf3), .Y(_311_) );
	AOI22X1 AOI22X1_22 ( .A(_1384_), .B(_1022__bF_buf2), .C(_268_), .D(_311_), .Y(_21_) );
	NAND3X1 NAND3X1_82 ( .A(_886__bF_buf3), .B(_1235_), .C(_280_), .Y(_312_) );
	OAI21X1 OAI21X1_258 ( .A(_1377_), .B(_886__bF_buf2), .C(_312_), .Y(_36_) );
	OAI21X1 OAI21X1_259 ( .A(_972_), .B(_1124_), .C(_882__bF_buf5), .Y(_313_) );
	NOR2X1 NOR2X1_164 ( .A(_881__bF_buf2), .B(_313_), .Y(_314_) );
	NAND2X1 NAND2X1_142 ( .A(D), .B(_1092_), .Y(_315_) );
	NOR2X1 NOR2X1_165 ( .A(_1203_), .B(_259_), .Y(_316_) );
	NAND2X1 NAND2X1_143 ( .A(_314_), .B(_316_), .Y(_317_) );
	OAI22X1 OAI22X1_32 ( .A(_152_), .B(_314_), .C(_315_), .D(_317_), .Y(_12_) );
	OAI21X1 OAI21X1_260 ( .A(_151_), .B(_314_), .C(_317_), .Y(_13_) );
	AOI22X1 AOI22X1_23 ( .A(_248_), .B(_305_), .C(_1100_), .D(_267_), .Y(_318_) );
	OAI21X1 OAI21X1_261 ( .A(_881__bF_buf1), .B(_885__bF_buf4), .C(inc), .Y(_319_) );
	OAI21X1 OAI21X1_262 ( .A(_1022__bF_buf1), .B(_318_), .C(_319_), .Y(_24_) );
	OAI21X1 OAI21X1_263 ( .A(_881__bF_buf0), .B(_885__bF_buf3), .C(load_only), .Y(_320_) );
	OAI21X1 OAI21X1_264 ( .A(_1022__bF_buf0), .B(_239_), .C(_320_), .Y(_26_) );
	INVX1 INVX1_104 ( .A(_1249_), .Y(_321_) );
	NAND3X1 NAND3X1_83 ( .A(_237_), .B(_1024_), .C(_321_), .Y(_322_) );
	OAI21X1 OAI21X1_265 ( .A(_986_), .B(_886__bF_buf1), .C(_322_), .Y(_40_) );
	NAND2X1 NAND2X1_144 ( .A(_177_), .B(_1466__bF_buf0), .Y(_323_) );
	NOR2X1 NOR2X1_166 ( .A(_1450_), .B(_323_), .Y(_324_) );
	NOR2X1 NOR2X1_167 ( .A(AXYS_1__0_), .B(_324_), .Y(_325_) );
	AOI21X1 AOI21X1_50 ( .A(_286_), .B(_324_), .C(_325_), .Y(_68_) );
	NAND2X1 NAND2X1_145 ( .A(_190_), .B(_324_), .Y(_326_) );
	OAI21X1 OAI21X1_266 ( .A(_1495_), .B(_324_), .C(_326_), .Y(_71_) );
	NOR2X1 NOR2X1_168 ( .A(AXYS_1__2_), .B(_324_), .Y(_327_) );
	AOI21X1 AOI21X1_51 ( .A(_292_), .B(_324_), .C(_327_), .Y(_74_) );
	NAND2X1 NAND2X1_146 ( .A(_324_), .B(_204_), .Y(_328_) );
	OAI21X1 OAI21X1_267 ( .A(_1520_), .B(_324_), .C(_328_), .Y(_76_) );
	NOR2X1 NOR2X1_169 ( .A(AXYS_1__4_), .B(_324_), .Y(_329_) );
	AOI21X1 AOI21X1_52 ( .A(_296_), .B(_324_), .C(_329_), .Y(_79_) );
	NOR2X1 NOR2X1_170 ( .A(AXYS_1__5_), .B(_324_), .Y(_330_) );
	AOI21X1 AOI21X1_53 ( .A(_217_), .B(_324_), .C(_330_), .Y(_82_) );
	NOR2X1 NOR2X1_171 ( .A(AXYS_1__6_), .B(_324_), .Y(_331_) );
	AOI21X1 AOI21X1_54 ( .A(_299_), .B(_324_), .C(_331_), .Y(_84_) );
	NAND2X1 NAND2X1_147 ( .A(_324_), .B(_229_), .Y(_332_) );
	OAI21X1 OAI21X1_268 ( .A(_72_), .B(_324_), .C(_332_), .Y(_86_) );
	NOR2X1 NOR2X1_172 ( .A(_1003_), .B(_237_), .Y(_333_) );
	OAI21X1 OAI21X1_269 ( .A(_919_), .B(_1148_), .C(_333_), .Y(_334_) );
	OAI21X1 OAI21X1_270 ( .A(_881__bF_buf7), .B(_885__bF_buf2), .C(store), .Y(_335_) );
	OAI21X1 OAI21X1_271 ( .A(_1022__bF_buf3), .B(_334_), .C(_335_), .Y(_39_) );
	OAI21X1 OAI21X1_272 ( .A(_881__bF_buf6), .B(_885__bF_buf1), .C(index_y), .Y(_336_) );
	OAI21X1 OAI21X1_273 ( .A(_1240_), .B(_1189_), .C(_886__bF_buf0), .Y(_337_) );
	NOR2X1 NOR2X1_173 ( .A(_237_), .B(_1249_), .Y(_338_) );
	NAND3X1 NAND3X1_84 ( .A(_898_), .B(_1024_), .C(_338_), .Y(_339_) );
	NAND3X1 NAND3X1_85 ( .A(_336_), .B(_339_), .C(_337_), .Y(_25_) );
	INVX1 INVX1_105 ( .A(src_reg_0_), .Y(_340_) );
	INVX1 INVX1_106 ( .A(_1254_), .Y(_341_) );
	NAND2X1 NAND2X1_148 ( .A(_924_), .B(_1100_), .Y(_342_) );
	OAI21X1 OAI21X1_274 ( .A(_910__bF_buf0), .B(_1002_), .C(_928_), .Y(_343_) );
	OR2X2 OR2X2_13 ( .A(_342_), .B(_343_), .Y(_344_) );
	OAI21X1 OAI21X1_275 ( .A(_1256_), .B(_264_), .C(_344_), .Y(_345_) );
	NAND2X1 NAND2X1_149 ( .A(_898_), .B(_333_), .Y(_346_) );
	INVX1 INVX1_107 ( .A(_270_), .Y(_347_) );
	NAND3X1 NAND3X1_86 ( .A(_995_), .B(_238_), .C(_347_), .Y(_348_) );
	OAI21X1 OAI21X1_276 ( .A(_1313_), .B(_346_), .C(_348_), .Y(_349_) );
	NOR2X1 NOR2X1_174 ( .A(_349_), .B(_345_), .Y(_350_) );
	OAI21X1 OAI21X1_277 ( .A(_341_), .B(_241_), .C(_350_), .Y(_351_) );
	NAND2X1 NAND2X1_150 ( .A(_886__bF_buf4), .B(_351_), .Y(_352_) );
	OAI21X1 OAI21X1_278 ( .A(_340_), .B(_886__bF_buf3), .C(_352_), .Y(_38__0_) );
	INVX1 INVX1_108 ( .A(src_reg_1_), .Y(_353_) );
	NAND2X1 NAND2X1_151 ( .A(_1257_), .B(_1254_), .Y(_354_) );
	OAI21X1 OAI21X1_279 ( .A(_266_), .B(_354_), .C(_886__bF_buf2), .Y(_355_) );
	NOR2X1 NOR2X1_175 ( .A(_1003_), .B(_904_), .Y(_356_) );
	OAI21X1 OAI21X1_280 ( .A(_347_), .B(_356_), .C(_338_), .Y(_357_) );
	OAI21X1 OAI21X1_281 ( .A(_1141_), .B(_264_), .C(_357_), .Y(_358_) );
	NOR2X1 NOR2X1_176 ( .A(_358_), .B(_355_), .Y(_359_) );
	AOI22X1 AOI22X1_24 ( .A(_353_), .B(_1022__bF_buf2), .C(_359_), .D(_350_), .Y(_38__1_) );
	INVX1 INVX1_109 ( .A(dst_reg_0_), .Y(_360_) );
	OAI21X1 OAI21X1_282 ( .A(_924_), .B(_908_), .C(_995_), .Y(_361_) );
	OAI21X1 OAI21X1_283 ( .A(_239_), .B(_361_), .C(_344_), .Y(_362_) );
	OAI21X1 OAI21X1_284 ( .A(_346_), .B(_341_), .C(_1230_), .Y(_363_) );
	OAI21X1 OAI21X1_285 ( .A(_363_), .B(_362_), .C(_886__bF_buf1), .Y(_364_) );
	OAI21X1 OAI21X1_286 ( .A(_360_), .B(_886__bF_buf0), .C(_364_), .Y(_23__0_) );
	INVX1 INVX1_110 ( .A(dst_reg_1_), .Y(_365_) );
	INVX1 INVX1_111 ( .A(_362_), .Y(_366_) );
	OAI22X1 OAI22X1_33 ( .A(_1249_), .B(_239_), .C(_1141_), .D(_249_), .Y(_367_) );
	NOR2X1 NOR2X1_177 ( .A(_355_), .B(_367_), .Y(_368_) );
	AOI22X1 AOI22X1_25 ( .A(_365_), .B(_1022__bF_buf1), .C(_368_), .D(_366_), .Y(_23__1_) );
	INVX1 INVX1_112 ( .A(load_reg), .Y(_369_) );
	NAND2X1 NAND2X1_152 ( .A(_1148_), .B(_240_), .Y(_370_) );
	NAND3X1 NAND3X1_87 ( .A(_1003_), .B(_1008_), .C(_930_), .Y(_371_) );
	OAI21X1 OAI21X1_287 ( .A(_910__bF_buf4), .B(_917_), .C(_1023_), .Y(_372_) );
	NOR2X1 NOR2X1_178 ( .A(_372_), .B(_237_), .Y(_373_) );
	AOI22X1 AOI22X1_26 ( .A(_356_), .B(_373_), .C(_999_), .D(_1254_), .Y(_374_) );
	NAND3X1 NAND3X1_88 ( .A(_371_), .B(_374_), .C(_370_), .Y(_375_) );
	NAND2X1 NAND2X1_153 ( .A(_1254_), .B(_240_), .Y(_376_) );
	NOR2X1 NOR2X1_179 ( .A(_1256_), .B(_266_), .Y(_377_) );
	AOI22X1 AOI22X1_27 ( .A(_919_), .B(_343_), .C(_1254_), .D(_377_), .Y(_378_) );
	NAND3X1 NAND3X1_89 ( .A(_342_), .B(_378_), .C(_376_), .Y(_379_) );
	OAI21X1 OAI21X1_288 ( .A(_375_), .B(_379_), .C(_886__bF_buf4), .Y(_380_) );
	OAI21X1 OAI21X1_289 ( .A(_369_), .B(_886__bF_buf3), .C(_380_), .Y(_27_) );
	NAND3X1 NAND3X1_90 ( .A(RDY_bF_buf5), .B(_1214_), .C(_1475_), .Y(_381_) );
	OAI21X1 OAI21X1_290 ( .A(_881__bF_buf5), .B(_885__bF_buf0), .C(IRHOLD_valid), .Y(_382_) );
	OAI21X1 OAI21X1_291 ( .A(reset), .B(_382_), .C(_381_), .Y(_5_) );
	NOR2X1 NOR2X1_180 ( .A(_1489_), .B(_323_), .Y(_383_) );
	NOR2X1 NOR2X1_181 ( .A(AXYS_3__0_), .B(_383_), .Y(_384_) );
	AOI21X1 AOI21X1_55 ( .A(_286_), .B(_383_), .C(_384_), .Y(_153_) );
	NOR2X1 NOR2X1_182 ( .A(AXYS_3__1_), .B(_383_), .Y(_385_) );
	AOI21X1 AOI21X1_56 ( .A(_290_), .B(_383_), .C(_385_), .Y(_154_) );
	NOR2X1 NOR2X1_183 ( .A(AXYS_3__2_), .B(_383_), .Y(_386_) );
	AOI21X1 AOI21X1_57 ( .A(_292_), .B(_383_), .C(_386_), .Y(_156_) );
	NOR2X1 NOR2X1_184 ( .A(AXYS_3__3_), .B(_383_), .Y(_387_) );
	AOI21X1 AOI21X1_58 ( .A(_294_), .B(_383_), .C(_387_), .Y(_159_) );
	NOR2X1 NOR2X1_185 ( .A(AXYS_3__4_), .B(_383_), .Y(_388_) );
	AOI21X1 AOI21X1_59 ( .A(_296_), .B(_383_), .C(_388_), .Y(_162_) );
	NOR2X1 NOR2X1_186 ( .A(AXYS_3__5_), .B(_383_), .Y(_389_) );
	AOI21X1 AOI21X1_60 ( .A(_217_), .B(_383_), .C(_389_), .Y(_165_) );
	NOR2X1 NOR2X1_187 ( .A(AXYS_3__6_), .B(_383_), .Y(_390_) );
	AOI21X1 AOI21X1_61 ( .A(_299_), .B(_383_), .C(_390_), .Y(_168_) );
	NOR2X1 NOR2X1_188 ( .A(AXYS_3__7_), .B(_383_), .Y(_391_) );
	AOI21X1 AOI21X1_62 ( .A(_301_), .B(_383_), .C(_391_), .Y(_171_) );
	NAND2X1 NAND2X1_154 ( .A(IRHOLD_0_), .B(_381_), .Y(_392_) );
	OAI21X1 OAI21X1_292 ( .A(_1403_), .B(_381_), .C(_392_), .Y(_4__0_) );
	NAND2X1 NAND2X1_155 ( .A(IRHOLD_1_), .B(_381_), .Y(_393_) );
	OAI21X1 OAI21X1_293 ( .A(_1419_), .B(_381_), .C(_393_), .Y(_4__1_) );
	NAND2X1 NAND2X1_156 ( .A(IRHOLD_2_), .B(_381_), .Y(_394_) );
	OAI21X1 OAI21X1_294 ( .A(_905_), .B(_381_), .C(_394_), .Y(_4__2_) );
	NAND2X1 NAND2X1_157 ( .A(IRHOLD_3_), .B(_381_), .Y(_395_) );
	OAI21X1 OAI21X1_295 ( .A(_1095_), .B(_381_), .C(_395_), .Y(_4__3_) );
	MUX2X1 MUX2X1_11 ( .A(_922_), .B(_891_), .S(_381_), .Y(_4__4_) );
	INVX1 INVX1_113 ( .A(IRHOLD_5_), .Y(_396_) );
	MUX2X1 MUX2X1_12 ( .A(_396_), .B(_1424_), .S(_381_), .Y(_4__5_) );
	MUX2X1 MUX2X1_13 ( .A(_1006_), .B(_1260_), .S(_381_), .Y(_4__6_) );
	INVX1 INVX1_114 ( .A(IRHOLD_7_), .Y(_397_) );
	MUX2X1 MUX2X1_14 ( .A(_397_), .B(_925_), .S(_381_), .Y(_4__7_) );
	NOR2X1 NOR2X1_189 ( .A(_255_), .B(_978_), .Y(_398_) );
	OAI21X1 OAI21X1_296 ( .A(_1038_), .B(_398_), .C(DIMUX_6_), .Y(_399_) );
	INVX1 INVX1_115 ( .A(_398_), .Y(_400_) );
	AOI21X1 AOI21X1_63 ( .A(_1177_), .B(_151_), .C(plp), .Y(_401_) );
	OAI21X1 OAI21X1_297 ( .A(_151_), .B(ALU_V), .C(_401_), .Y(_402_) );
	OAI22X1 OAI22X1_34 ( .A(_224_), .B(_158_), .C(clv), .D(_402_), .Y(_403_) );
	NOR2X1 NOR2X1_190 ( .A(_1177_), .B(_1436_), .Y(_404_) );
	AOI22X1 AOI22X1_28 ( .A(_1436_), .B(_403_), .C(_404_), .D(_400_), .Y(_405_) );
	OAI21X1 OAI21X1_298 ( .A(_1038_), .B(_405_), .C(_399_), .Y(_10_) );
	NOR2X1 NOR2X1_191 ( .A(plp), .B(cld), .Y(_406_) );
	OAI21X1 OAI21X1_299 ( .A(D), .B(sed), .C(_406_), .Y(_407_) );
	OAI21X1 OAI21X1_300 ( .A(_199_), .B(_158_), .C(_407_), .Y(_408_) );
	OAI21X1 OAI21X1_301 ( .A(_124_), .B(_1436_), .C(_1392_), .Y(_409_) );
	AOI21X1 AOI21X1_64 ( .A(_1436_), .B(_408_), .C(_409_), .Y(_410_) );
	AOI21X1 AOI21X1_65 ( .A(_1095_), .B(_1038_), .C(_410_), .Y(_3_) );
	NAND2X1 NAND2X1_158 ( .A(ALU_N), .B(_959_), .Y(_411_) );
	INVX1 INVX1_116 ( .A(_1449_), .Y(_412_) );
	NAND2X1 NAND2X1_159 ( .A(_412_), .B(_1459_), .Y(_413_) );
	NAND3X1 NAND3X1_91 ( .A(_1440_), .B(_413_), .C(_1466__bF_buf4), .Y(_414_) );
	AOI21X1 AOI21X1_66 ( .A(_414_), .B(load_reg), .C(compare), .Y(_415_) );
	NAND2X1 NAND2X1_160 ( .A(N), .B(_415_), .Y(_416_) );
	OAI21X1 OAI21X1_302 ( .A(_1450_), .B(_1470_), .C(load_reg), .Y(_417_) );
	NAND2X1 NAND2X1_161 ( .A(_1384_), .B(_417_), .Y(_418_) );
	AOI21X1 AOI21X1_67 ( .A(_418_), .B(ALU_N), .C(plp), .Y(_419_) );
	NAND2X1 NAND2X1_162 ( .A(_416_), .B(_419_), .Y(_420_) );
	INVX1 INVX1_117 ( .A(ADD_7_), .Y(_421_) );
	AOI21X1 AOI21X1_68 ( .A(_421_), .B(plp), .C(_885__bF_buf4), .Y(_422_) );
	NAND2X1 NAND2X1_163 ( .A(_925_), .B(_398_), .Y(_423_) );
	OAI21X1 OAI21X1_303 ( .A(N), .B(_398_), .C(_423_), .Y(_424_) );
	OAI21X1 OAI21X1_304 ( .A(_1436_), .B(_424_), .C(_1392_), .Y(_425_) );
	AOI21X1 AOI21X1_69 ( .A(_420_), .B(_422_), .C(_425_), .Y(_426_) );
	OAI21X1 OAI21X1_305 ( .A(DIMUX_7_), .B(_1392_), .C(_95_), .Y(_427_) );
	OAI21X1 OAI21X1_306 ( .A(_427_), .B(_426_), .C(_411_), .Y(_8_) );
	NAND2X1 NAND2X1_164 ( .A(ALU_Z), .B(_959_), .Y(_428_) );
	NAND3X1 NAND3X1_92 ( .A(_1384_), .B(_255_), .C(_417_), .Y(_429_) );
	NAND2X1 NAND2X1_165 ( .A(ALU_Z), .B(_429_), .Y(_430_) );
	NAND3X1 NAND3X1_93 ( .A(Z), .B(_255_), .C(_415_), .Y(_431_) );
	NAND3X1 NAND3X1_94 ( .A(_158_), .B(_430_), .C(_431_), .Y(_432_) );
	INVX2 INVX2_37 ( .A(ADD_1_), .Y(_433_) );
	AOI21X1 AOI21X1_70 ( .A(_433_), .B(plp), .C(_885__bF_buf3), .Y(_434_) );
	OAI21X1 OAI21X1_307 ( .A(_1174_), .B(_1436_), .C(_1392_), .Y(_435_) );
	AOI21X1 AOI21X1_71 ( .A(_432_), .B(_434_), .C(_435_), .Y(_436_) );
	OAI21X1 OAI21X1_308 ( .A(DIMUX_1_), .B(_1392_), .C(_95_), .Y(_437_) );
	OAI21X1 OAI21X1_309 ( .A(_437_), .B(_436_), .C(_428_), .Y(_11_) );
	INVX1 INVX1_118 ( .A(ALU_CO), .Y(_438_) );
	NAND2X1 NAND2X1_166 ( .A(shift), .B(_959_), .Y(_439_) );
	NOR2X1 NOR2X1_192 ( .A(write_back), .B(_885__bF_buf2), .Y(_440_) );
	NAND3X1 NAND3X1_95 ( .A(_1377_), .B(_1384_), .C(_151_), .Y(_441_) );
	NAND2X1 NAND2X1_167 ( .A(_1376_), .B(_251_), .Y(_442_) );
	NOR2X1 NOR2X1_193 ( .A(plp), .B(clc), .Y(_443_) );
	AOI22X1 AOI22X1_29 ( .A(ADD_0_), .B(plp), .C(_443_), .D(_442_), .Y(_444_) );
	NAND2X1 NAND2X1_168 ( .A(ALU_CO), .B(_441_), .Y(_445_) );
	OAI21X1 OAI21X1_310 ( .A(_441_), .B(_444_), .C(_445_), .Y(_446_) );
	OAI21X1 OAI21X1_311 ( .A(_1376_), .B(_440_), .C(_1392_), .Y(_447_) );
	AOI21X1 AOI21X1_72 ( .A(_446_), .B(_440_), .C(_447_), .Y(_448_) );
	OAI21X1 OAI21X1_312 ( .A(DIMUX_0_), .B(_1392_), .C(_439_), .Y(_449_) );
	OAI22X1 OAI22X1_35 ( .A(_438_), .B(_439_), .C(_449_), .D(_448_), .Y(_2_) );
	NAND2X1 NAND2X1_169 ( .A(RDY_bF_buf4), .B(DI[7]), .Y(_450_) );
	OAI21X1 OAI21X1_313 ( .A(RDY_bF_buf3), .B(_85_), .C(_450_), .Y(_15_) );
	OAI21X1 OAI21X1_314 ( .A(_1027_), .B(_962__bF_buf1), .C(_1392_), .Y(_451_) );
	AOI21X1 AOI21X1_73 ( .A(_963_), .B(_1043_), .C(_451_), .Y(_452_) );
	NAND3X1 NAND3X1_96 ( .A(_1429_), .B(_1457_), .C(_452_), .Y(_453_) );
	OAI21X1 OAI21X1_315 ( .A(_947_), .B(_956_), .C(_1192_), .Y(_454_) );
	OAI21X1 OAI21X1_316 ( .A(state_5_), .B(_936__bF_buf1), .C(_454_), .Y(_455_) );
	AOI21X1 AOI21X1_74 ( .A(_882__bF_buf4), .B(_984_), .C(_1032_), .Y(_456_) );
	OAI21X1 OAI21X1_317 ( .A(_1209_), .B(_962__bF_buf0), .C(_456_), .Y(_457_) );
	NOR2X1 NOR2X1_194 ( .A(_455_), .B(_457_), .Y(_458_) );
	NOR2X1 NOR2X1_195 ( .A(_1075_), .B(_1028_), .Y(_459_) );
	OAI21X1 OAI21X1_318 ( .A(_936__bF_buf0), .B(_945_), .C(_459_), .Y(_460_) );
	NOR2X1 NOR2X1_196 ( .A(_1112_), .B(_460_), .Y(_461_) );
	NAND2X1 NAND2X1_170 ( .A(_461_), .B(_458_), .Y(_462_) );
	NOR2X1 NOR2X1_197 ( .A(_453_), .B(_462_), .Y(_463_) );
	OAI21X1 OAI21X1_319 ( .A(_957__bF_buf4), .B(_958_), .C(_1378_), .Y(_464_) );
	OR2X2 OR2X2_14 ( .A(_464_), .B(_1224_), .Y(_465_) );
	NOR2X1 NOR2X1_198 ( .A(_1397_), .B(_87_), .Y(_466_) );
	NOR2X1 NOR2X1_199 ( .A(_1068_), .B(_967_), .Y(_467_) );
	OAI21X1 OAI21X1_320 ( .A(_937__bF_buf2), .B(_1209_), .C(_467_), .Y(_468_) );
	OAI21X1 OAI21X1_321 ( .A(_962__bF_buf4), .B(_1076_), .C(_951_), .Y(_469_) );
	NOR2X1 NOR2X1_200 ( .A(_469_), .B(_468_), .Y(_470_) );
	NAND2X1 NAND2X1_171 ( .A(_466_), .B(_470_), .Y(_471_) );
	NOR2X1 NOR2X1_201 ( .A(_465_), .B(_471_), .Y(_472_) );
	NAND2X1 NAND2X1_172 ( .A(_463_), .B(_472_), .Y(_473_) );
	INVX2 INVX2_38 ( .A(_458_), .Y(_474_) );
	AOI22X1 AOI22X1_30 ( .A(_464_), .B(ABH_0_), .C(ADD_0_), .D(_468_), .Y(_475_) );
	NAND3X1 NAND3X1_97 ( .A(_1433_), .B(_466_), .C(_475_), .Y(_476_) );
	OR2X2 OR2X2_15 ( .A(_476_), .B(_453_), .Y(_477_) );
	AOI21X1 AOI21X1_75 ( .A(DIMUX_0_), .B(_474_), .C(_477_), .Y(_478_) );
	OAI21X1 OAI21X1_322 ( .A(_102_), .B(_473_), .C(_478_), .Y(_1536__8_) );
	INVX1 INVX1_119 ( .A(ABH_0_), .Y(_479_) );
	OAI21X1 OAI21X1_323 ( .A(_961_), .B(_1043_), .C(_963_), .Y(_480_) );
	NAND3X1 NAND3X1_98 ( .A(_480_), .B(_456_), .C(_467_), .Y(_481_) );
	NOR2X1 NOR2X1_202 ( .A(_1073_), .B(_977_), .Y(_482_) );
	NOR3X1 NOR3X1_16 ( .A(state_3_), .B(_964_), .C(_949_), .Y(_483_) );
	OAI21X1 OAI21X1_324 ( .A(_950_), .B(_483_), .C(_947_), .Y(_484_) );
	NAND2X1 NAND2X1_173 ( .A(_484_), .B(_482_), .Y(_485_) );
	INVX1 INVX1_120 ( .A(_485_), .Y(_486_) );
	NAND3X1 NAND3X1_99 ( .A(_1456_), .B(_459_), .C(_486_), .Y(_487_) );
	NOR2X1 NOR2X1_203 ( .A(_481_), .B(_487_), .Y(_488_) );
	NOR2X1 NOR2X1_204 ( .A(_1198_), .B(_1194_), .Y(_489_) );
	AOI21X1 AOI21X1_76 ( .A(_946_), .B(_1215_), .C(_1128_), .Y(_490_) );
	NAND3X1 NAND3X1_100 ( .A(_490_), .B(_489_), .C(_1220_), .Y(_491_) );
	NOR2X1 NOR2X1_205 ( .A(_1108_), .B(_1120_), .Y(_492_) );
	NOR2X1 NOR2X1_206 ( .A(_1112_), .B(_1282_), .Y(_493_) );
	NAND2X1 NAND2X1_174 ( .A(_492_), .B(_493_), .Y(_494_) );
	AOI21X1 AOI21X1_77 ( .A(_945_), .B(_972_), .C(_1388_), .Y(_495_) );
	OAI21X1 OAI21X1_325 ( .A(state_5_), .B(_1119_), .C(_495_), .Y(_496_) );
	OR2X2 OR2X2_16 ( .A(_496_), .B(_494_), .Y(_497_) );
	NOR2X1 NOR2X1_207 ( .A(_491_), .B(_497_), .Y(_498_) );
	AOI22X1 AOI22X1_31 ( .A(_955_), .B(_1453_), .C(_956_), .D(_1034__bF_buf3), .Y(_499_) );
	OAI21X1 OAI21X1_326 ( .A(_936__bF_buf3), .B(_937__bF_buf1), .C(_499_), .Y(_500_) );
	OAI21X1 OAI21X1_327 ( .A(state_4_), .B(_966_), .C(_454_), .Y(_501_) );
	OAI21X1 OAI21X1_328 ( .A(_936__bF_buf2), .B(_882__bF_buf3), .C(_1193_), .Y(_502_) );
	NOR2X1 NOR2X1_208 ( .A(_502_), .B(_501_), .Y(_503_) );
	AOI22X1 AOI22X1_32 ( .A(_1034__bF_buf2), .B(_955_), .C(_963_), .D(_1046_), .Y(_504_) );
	NAND2X1 NAND2X1_175 ( .A(_504_), .B(_503_), .Y(_505_) );
	NOR2X1 NOR2X1_209 ( .A(_500_), .B(_505_), .Y(_506_) );
	NAND3X1 NAND3X1_101 ( .A(_1080_), .B(_499_), .C(_504_), .Y(_507_) );
	OAI21X1 OAI21X1_329 ( .A(_936__bF_buf1), .B(_947_), .C(_1193_), .Y(_508_) );
	OR2X2 OR2X2_17 ( .A(_501_), .B(_508_), .Y(_509_) );
	NOR2X1 NOR2X1_210 ( .A(_507_), .B(_509_), .Y(_510_) );
	OAI21X1 OAI21X1_330 ( .A(_510_), .B(_506_), .C(_498_), .Y(_511_) );
	OAI21X1 OAI21X1_331 ( .A(_957__bF_buf3), .B(_1111_), .C(_490_), .Y(_512_) );
	INVX1 INVX1_121 ( .A(_1188_), .Y(_513_) );
	NOR2X1 NOR2X1_211 ( .A(_1128_), .B(_1388_), .Y(_514_) );
	NAND3X1 NAND3X1_102 ( .A(_513_), .B(_313_), .C(_514_), .Y(_515_) );
	INVX1 INVX1_122 ( .A(_1271_), .Y(_516_) );
	NOR2X1 NOR2X1_212 ( .A(_1132_), .B(_1198_), .Y(_517_) );
	NAND3X1 NAND3X1_103 ( .A(_516_), .B(_1483_), .C(_517_), .Y(_518_) );
	OAI22X1 OAI22X1_36 ( .A(_496_), .B(_512_), .C(_518_), .D(_515_), .Y(_519_) );
	NOR2X1 NOR2X1_213 ( .A(_1219_), .B(_1407_), .Y(_520_) );
	NAND3X1 NAND3X1_104 ( .A(_1396_), .B(_1405_), .C(_520_), .Y(_521_) );
	OR2X2 OR2X2_18 ( .A(_494_), .B(_500_), .Y(_522_) );
	NOR2X1 NOR2X1_214 ( .A(_521_), .B(_522_), .Y(_523_) );
	NAND3X1 NAND3X1_105 ( .A(_503_), .B(_519_), .C(_523_), .Y(_524_) );
	NAND2X1 NAND2X1_176 ( .A(_524_), .B(_511_), .Y(_525_) );
	OR2X2 OR2X2_19 ( .A(_481_), .B(_485_), .Y(_526_) );
	OR2X2 OR2X2_20 ( .A(_526_), .B(_507_), .Y(_527_) );
	OAI21X1 OAI21X1_332 ( .A(_936__bF_buf0), .B(_957__bF_buf2), .C(_1193_), .Y(_528_) );
	OAI21X1 OAI21X1_333 ( .A(state_5_), .B(_936__bF_buf3), .C(_1053_), .Y(_529_) );
	OR2X2 OR2X2_21 ( .A(_529_), .B(_528_), .Y(_530_) );
	OR2X2 OR2X2_22 ( .A(_530_), .B(_460_), .Y(_531_) );
	NOR2X1 NOR2X1_215 ( .A(_501_), .B(_531_), .Y(_532_) );
	NAND2X1 NAND2X1_177 ( .A(_498_), .B(_532_), .Y(_533_) );
	OAI21X1 OAI21X1_334 ( .A(_527_), .B(_533_), .C(RDY_bF_buf2), .Y(_534_) );
	AOI21X1 AOI21X1_78 ( .A(_525_), .B(_488_), .C(_534_), .Y(_535_) );
	NAND2X1 NAND2X1_178 ( .A(_1536__8_), .B(_535__bF_buf4), .Y(_536_) );
	OAI21X1 OAI21X1_335 ( .A(_479_), .B(_535__bF_buf3), .C(_536_), .Y(_0__0_) );
	INVX4 INVX4_14 ( .A(_468_), .Y(_537_) );
	OAI21X1 OAI21X1_336 ( .A(_1224_), .B(_464_), .C(ABH_1_), .Y(_538_) );
	OAI21X1 OAI21X1_337 ( .A(_433_), .B(_537_), .C(_538_), .Y(_539_) );
	AOI21X1 AOI21X1_79 ( .A(DIMUX_1_), .B(_474_), .C(_539_), .Y(_540_) );
	OAI21X1 OAI21X1_338 ( .A(_107_), .B(_473_), .C(_540_), .Y(_1536__9_) );
	INVX1 INVX1_123 ( .A(ABH_1_), .Y(_541_) );
	NAND2X1 NAND2X1_179 ( .A(_1536__9_), .B(_535__bF_buf2), .Y(_542_) );
	OAI21X1 OAI21X1_339 ( .A(_541_), .B(_535__bF_buf1), .C(_542_), .Y(_0__1_) );
	OAI22X1 OAI22X1_37 ( .A(_115_), .B(_537_), .C(_905_), .D(_458_), .Y(_543_) );
	AOI21X1 AOI21X1_80 ( .A(ABH_2_), .B(_465_), .C(_543_), .Y(_544_) );
	OAI21X1 OAI21X1_340 ( .A(_114_), .B(_473_), .C(_544_), .Y(_1536__10_) );
	INVX1 INVX1_124 ( .A(ABH_2_), .Y(_545_) );
	NAND2X1 NAND2X1_180 ( .A(_1536__10_), .B(_535__bF_buf0), .Y(_546_) );
	OAI21X1 OAI21X1_341 ( .A(_545_), .B(_535__bF_buf4), .C(_546_), .Y(_0__2_) );
	OAI22X1 OAI22X1_38 ( .A(_199_), .B(_537_), .C(_1095_), .D(_458_), .Y(_547_) );
	AOI21X1 AOI21X1_81 ( .A(ABH_3_), .B(_465_), .C(_547_), .Y(_548_) );
	OAI21X1 OAI21X1_342 ( .A(_122_), .B(_473_), .C(_548_), .Y(_1536__11_) );
	INVX1 INVX1_125 ( .A(ABH_3_), .Y(_549_) );
	NAND2X1 NAND2X1_181 ( .A(_1536__11_), .B(_535__bF_buf3), .Y(_550_) );
	OAI21X1 OAI21X1_343 ( .A(_549_), .B(_535__bF_buf2), .C(_550_), .Y(_0__3_) );
	INVX1 INVX1_126 ( .A(ADD_4_), .Y(_551_) );
	OAI22X1 OAI22X1_39 ( .A(_551_), .B(_537_), .C(_891_), .D(_458_), .Y(_552_) );
	AOI21X1 AOI21X1_82 ( .A(ABH_4_), .B(_465_), .C(_552_), .Y(_553_) );
	OAI21X1 OAI21X1_344 ( .A(_131_), .B(_473_), .C(_553_), .Y(_1536__12_) );
	NAND2X1 NAND2X1_182 ( .A(_1536__12_), .B(_535__bF_buf1), .Y(_554_) );
	OAI21X1 OAI21X1_345 ( .A(_1525_), .B(_535__bF_buf0), .C(_554_), .Y(_0__4_) );
	OAI21X1 OAI21X1_346 ( .A(_1224_), .B(_464_), .C(ABH_5_), .Y(_555_) );
	OAI21X1 OAI21X1_347 ( .A(_209_), .B(_537_), .C(_555_), .Y(_556_) );
	AOI21X1 AOI21X1_83 ( .A(DIMUX_5_), .B(_474_), .C(_556_), .Y(_557_) );
	OAI21X1 OAI21X1_348 ( .A(_135_), .B(_473_), .C(_557_), .Y(_1536__13_) );
	NAND2X1 NAND2X1_183 ( .A(_1536__13_), .B(_535__bF_buf4), .Y(_558_) );
	OAI21X1 OAI21X1_349 ( .A(_42_), .B(_535__bF_buf3), .C(_558_), .Y(_0__5_) );
	OAI22X1 OAI22X1_40 ( .A(_224_), .B(_537_), .C(_1260_), .D(_458_), .Y(_559_) );
	AOI21X1 AOI21X1_84 ( .A(ABH_6_), .B(_465_), .C(_559_), .Y(_560_) );
	OAI21X1 OAI21X1_350 ( .A(_142_), .B(_473_), .C(_560_), .Y(_1536__14_) );
	NAND2X1 NAND2X1_184 ( .A(_1536__14_), .B(_535__bF_buf2), .Y(_561_) );
	OAI21X1 OAI21X1_351 ( .A(_52_), .B(_535__bF_buf1), .C(_561_), .Y(_0__6_) );
	OAI21X1 OAI21X1_352 ( .A(_1224_), .B(_464_), .C(ABH_7_), .Y(_562_) );
	OAI21X1 OAI21X1_353 ( .A(_421_), .B(_537_), .C(_562_), .Y(_563_) );
	AOI21X1 AOI21X1_85 ( .A(DIMUX_7_), .B(_474_), .C(_563_), .Y(_564_) );
	OAI21X1 OAI21X1_354 ( .A(_147_), .B(_473_), .C(_564_), .Y(_1536__15_) );
	NAND2X1 NAND2X1_185 ( .A(_1536__15_), .B(_535__bF_buf0), .Y(_565_) );
	OAI21X1 OAI21X1_355 ( .A(_62_), .B(_535__bF_buf4), .C(_565_), .Y(_0__7_) );
	NOR2X1 NOR2X1_216 ( .A(_466_), .B(_1474_), .Y(_566_) );
	INVX4 INVX4_15 ( .A(_463_), .Y(_567_) );
	INVX1 INVX1_127 ( .A(ABL_0_), .Y(_568_) );
	AOI22X1 AOI22X1_33 ( .A(ADD_0_), .B(_1224_), .C(DIMUX_0_), .D(_469_), .Y(_569_) );
	NOR2X1 NOR2X1_217 ( .A(_464_), .B(_468_), .Y(_570_) );
	OAI21X1 OAI21X1_356 ( .A(_568_), .B(_570_), .C(_569_), .Y(_571_) );
	AOI21X1 AOI21X1_86 ( .A(_567_), .B(ADD_0_), .C(_571_), .Y(_572_) );
	OAI21X1 OAI21X1_357 ( .A(_1402_), .B(_473_), .C(_572_), .Y(_573_) );
	OR2X2 OR2X2_23 ( .A(_573_), .B(_566_), .Y(_1536__0_) );
	OAI21X1 OAI21X1_358 ( .A(_566_), .B(_573_), .C(_535__bF_buf3), .Y(_574_) );
	OAI21X1 OAI21X1_359 ( .A(_568_), .B(_535__bF_buf2), .C(_574_), .Y(_1__0_) );
	NOR2X1 NOR2X1_218 ( .A(_466_), .B(_1497_), .Y(_575_) );
	INVX1 INVX1_128 ( .A(ABL_1_), .Y(_576_) );
	AOI22X1 AOI22X1_34 ( .A(_1224_), .B(ADD_1_), .C(DIMUX_1_), .D(_469_), .Y(_577_) );
	OAI21X1 OAI21X1_360 ( .A(_576_), .B(_570_), .C(_577_), .Y(_578_) );
	AOI21X1 AOI21X1_87 ( .A(_567_), .B(ADD_1_), .C(_578_), .Y(_579_) );
	OAI21X1 OAI21X1_361 ( .A(_1418_), .B(_473_), .C(_579_), .Y(_580_) );
	OR2X2 OR2X2_24 ( .A(_580_), .B(_575_), .Y(_1536__1_) );
	OAI21X1 OAI21X1_362 ( .A(_575_), .B(_580_), .C(_535__bF_buf1), .Y(_581_) );
	OAI21X1 OAI21X1_363 ( .A(_576_), .B(_535__bF_buf0), .C(_581_), .Y(_1__1_) );
	NOR2X1 NOR2X1_219 ( .A(_466_), .B(_1507_), .Y(_582_) );
	INVX1 INVX1_129 ( .A(ABL_2_), .Y(_583_) );
	AOI22X1 AOI22X1_35 ( .A(_1224_), .B(ADD_2_), .C(DIMUX_2_), .D(_469_), .Y(_584_) );
	OAI21X1 OAI21X1_364 ( .A(_583_), .B(_570_), .C(_584_), .Y(_585_) );
	AOI21X1 AOI21X1_88 ( .A(_567_), .B(ADD_2_), .C(_585_), .Y(_586_) );
	OAI21X1 OAI21X1_365 ( .A(_1420_), .B(_473_), .C(_586_), .Y(_587_) );
	OR2X2 OR2X2_25 ( .A(_587_), .B(_582_), .Y(_1536__2_) );
	OAI21X1 OAI21X1_366 ( .A(_582_), .B(_587_), .C(_535__bF_buf4), .Y(_588_) );
	OAI21X1 OAI21X1_367 ( .A(_583_), .B(_535__bF_buf3), .C(_588_), .Y(_1__2_) );
	NOR2X1 NOR2X1_220 ( .A(_466_), .B(_1523_), .Y(_589_) );
	INVX1 INVX1_130 ( .A(ABL_3_), .Y(_590_) );
	AOI22X1 AOI22X1_36 ( .A(_1224_), .B(ADD_3_), .C(DIMUX_3_), .D(_469_), .Y(_591_) );
	OAI21X1 OAI21X1_368 ( .A(_590_), .B(_570_), .C(_591_), .Y(_592_) );
	AOI21X1 AOI21X1_89 ( .A(_567_), .B(ADD_3_), .C(_592_), .Y(_593_) );
	OAI21X1 OAI21X1_369 ( .A(_1421_), .B(_473_), .C(_593_), .Y(_594_) );
	OR2X2 OR2X2_26 ( .A(_594_), .B(_589_), .Y(_1536__3_) );
	OAI21X1 OAI21X1_370 ( .A(_589_), .B(_594_), .C(_535__bF_buf2), .Y(_595_) );
	OAI21X1 OAI21X1_371 ( .A(_590_), .B(_535__bF_buf1), .C(_595_), .Y(_1__3_) );
	NOR2X1 NOR2X1_221 ( .A(_466_), .B(_41_), .Y(_596_) );
	INVX1 INVX1_131 ( .A(ABL_4_), .Y(_597_) );
	AOI22X1 AOI22X1_37 ( .A(_1224_), .B(ADD_4_), .C(DIMUX_4_), .D(_469_), .Y(_598_) );
	OAI21X1 OAI21X1_372 ( .A(_597_), .B(_570_), .C(_598_), .Y(_599_) );
	AOI21X1 AOI21X1_90 ( .A(_567_), .B(ADD_4_), .C(_599_), .Y(_600_) );
	OAI21X1 OAI21X1_373 ( .A(_1422_), .B(_473_), .C(_600_), .Y(_601_) );
	OR2X2 OR2X2_27 ( .A(_601_), .B(_596_), .Y(_1536__4_) );
	OAI21X1 OAI21X1_374 ( .A(_596_), .B(_601_), .C(_535__bF_buf0), .Y(_602_) );
	OAI21X1 OAI21X1_375 ( .A(_597_), .B(_535__bF_buf4), .C(_602_), .Y(_1__4_) );
	NOR2X1 NOR2X1_222 ( .A(_466_), .B(_51_), .Y(_603_) );
	INVX1 INVX1_132 ( .A(ABL_5_), .Y(_604_) );
	AOI22X1 AOI22X1_38 ( .A(_1224_), .B(ADD_5_), .C(DIMUX_5_), .D(_469_), .Y(_605_) );
	OAI21X1 OAI21X1_376 ( .A(_604_), .B(_570_), .C(_605_), .Y(_606_) );
	AOI21X1 AOI21X1_91 ( .A(_567_), .B(ADD_5_), .C(_606_), .Y(_607_) );
	OAI21X1 OAI21X1_377 ( .A(_1423_), .B(_473_), .C(_607_), .Y(_608_) );
	OR2X2 OR2X2_28 ( .A(_608_), .B(_603_), .Y(_1536__5_) );
	OAI21X1 OAI21X1_378 ( .A(_603_), .B(_608_), .C(_535__bF_buf3), .Y(_609_) );
	OAI21X1 OAI21X1_379 ( .A(_604_), .B(_535__bF_buf2), .C(_609_), .Y(_1__5_) );
	NOR2X1 NOR2X1_223 ( .A(_466_), .B(_61_), .Y(_610_) );
	INVX1 INVX1_133 ( .A(ABL_6_), .Y(_611_) );
	AOI22X1 AOI22X1_39 ( .A(_1224_), .B(ADD_6_), .C(DIMUX_6_), .D(_469_), .Y(_612_) );
	OAI21X1 OAI21X1_380 ( .A(_611_), .B(_570_), .C(_612_), .Y(_613_) );
	AOI21X1 AOI21X1_92 ( .A(_567_), .B(ADD_6_), .C(_613_), .Y(_614_) );
	OAI21X1 OAI21X1_381 ( .A(_1425_), .B(_473_), .C(_614_), .Y(_615_) );
	OR2X2 OR2X2_29 ( .A(_615_), .B(_610_), .Y(_1536__6_) );
	OAI21X1 OAI21X1_382 ( .A(_610_), .B(_615_), .C(_535__bF_buf1), .Y(_616_) );
	OAI21X1 OAI21X1_383 ( .A(_611_), .B(_535__bF_buf0), .C(_616_), .Y(_1__6_) );
	NOR2X1 NOR2X1_224 ( .A(_466_), .B(_75_), .Y(_617_) );
	INVX1 INVX1_134 ( .A(ABL_7_), .Y(_618_) );
	AOI22X1 AOI22X1_40 ( .A(_1224_), .B(ADD_7_), .C(DIMUX_7_), .D(_469_), .Y(_619_) );
	OAI21X1 OAI21X1_384 ( .A(_618_), .B(_570_), .C(_619_), .Y(_620_) );
	AOI21X1 AOI21X1_93 ( .A(_567_), .B(ADD_7_), .C(_620_), .Y(_621_) );
	OAI21X1 OAI21X1_385 ( .A(_1426_), .B(_473_), .C(_621_), .Y(_622_) );
	OR2X2 OR2X2_30 ( .A(_622_), .B(_617_), .Y(_1536__7_) );
	OAI21X1 OAI21X1_386 ( .A(_617_), .B(_622_), .C(_535__bF_buf4), .Y(_623_) );
	OAI21X1 OAI21X1_387 ( .A(_618_), .B(_535__bF_buf3), .C(_623_), .Y(_1__7_) );
	AND2X2 AND2X2_34 ( .A(_957__bF_buf1), .B(_962__bF_buf3), .Y(_624_) );
	NOR2X1 NOR2X1_225 ( .A(_1117_), .B(_624_), .Y(_625_) );
	OAI22X1 OAI22X1_41 ( .A(_962__bF_buf2), .B(_1031_), .C(_971_), .D(_624_), .Y(_626_) );
	NOR2X1 NOR2X1_226 ( .A(_625_), .B(_626_), .Y(_627_) );
	OAI21X1 OAI21X1_388 ( .A(_972_), .B(_1046_), .C(_882__bF_buf2), .Y(_628_) );
	OAI21X1 OAI21X1_389 ( .A(_483_), .B(_1034__bF_buf1), .C(_882__bF_buf1), .Y(_629_) );
	AND2X2 AND2X2_35 ( .A(_628_), .B(_629_), .Y(_630_) );
	NAND2X1 NAND2X1_186 ( .A(_627_), .B(_630_), .Y(_631_) );
	AOI22X1 AOI22X1_41 ( .A(_483_), .B(_956_), .C(_961_), .D(_963_), .Y(_632_) );
	OAI21X1 OAI21X1_390 ( .A(_624_), .B(_1117_), .C(_632_), .Y(_633_) );
	NAND3X1 NAND3X1_106 ( .A(ADD_0_), .B(_882__bF_buf0), .C(_1034__bF_buf0), .Y(_634_) );
	NAND3X1 NAND3X1_107 ( .A(PC_0_), .B(_882__bF_buf5), .C(_483_), .Y(_635_) );
	NAND2X1 NAND2X1_187 ( .A(ABL_0_), .B(_910__bF_buf3), .Y(_636_) );
	OAI21X1 OAI21X1_391 ( .A(_1402_), .B(_910__bF_buf2), .C(_636_), .Y(_637_) );
	NAND2X1 NAND2X1_188 ( .A(_1436_), .B(_637_), .Y(_638_) );
	NAND3X1 NAND3X1_108 ( .A(_634_), .B(_635_), .C(_638_), .Y(_639_) );
	AOI21X1 AOI21X1_94 ( .A(ADD_0_), .B(_633_), .C(_639_), .Y(_640_) );
	OAI21X1 OAI21X1_392 ( .A(_1402_), .B(_631_), .C(_640_), .Y(_641_) );
	NOR2X1 NOR2X1_227 ( .A(_910__bF_buf1), .B(_885__bF_buf1), .Y(_642_) );
	OAI21X1 OAI21X1_393 ( .A(_1064_), .B(_1065_), .C(_454_), .Y(_643_) );
	NOR2X1 NOR2X1_228 ( .A(_642_), .B(_643_), .Y(_644_) );
	OAI21X1 OAI21X1_394 ( .A(_937__bF_buf0), .B(_1051_), .C(_1127_), .Y(_645_) );
	OAI22X1 OAI22X1_42 ( .A(state_5_), .B(_1031_), .C(state_4_), .D(_971_), .Y(_646_) );
	NOR2X1 NOR2X1_229 ( .A(_645_), .B(_646_), .Y(_647_) );
	OAI21X1 OAI21X1_395 ( .A(_937__bF_buf4), .B(_1076_), .C(_1103_), .Y(_648_) );
	INVX1 INVX1_135 ( .A(_648_), .Y(_649_) );
	NAND3X1 NAND3X1_109 ( .A(_647_), .B(_649_), .C(_644_), .Y(_650_) );
	NOR2X1 NOR2X1_230 ( .A(_650_), .B(_641_), .Y(_651_) );
	NAND2X1 NAND2X1_189 ( .A(_628_), .B(_629_), .Y(_652_) );
	NOR3X1 NOR3X1_17 ( .A(_1402_), .B(_633_), .C(_652_), .Y(_653_) );
	OAI21X1 OAI21X1_396 ( .A(_625_), .B(_626_), .C(ADD_0_), .Y(_654_) );
	AND2X2 AND2X2_36 ( .A(_634_), .B(_635_), .Y(_655_) );
	NAND3X1 NAND3X1_110 ( .A(_638_), .B(_655_), .C(_654_), .Y(_656_) );
	OAI21X1 OAI21X1_397 ( .A(_656_), .B(_653_), .C(_650_), .Y(_657_) );
	NAND2X1 NAND2X1_190 ( .A(RDY_bF_buf1), .B(_657_), .Y(_658_) );
	OAI22X1 OAI22X1_43 ( .A(RDY_bF_buf0), .B(_1402_), .C(_658_), .D(_651_), .Y(_9__0_) );
	NAND3X1 NAND3X1_111 ( .A(PC_0_), .B(_627_), .C(_630_), .Y(_659_) );
	AND2X2 AND2X2_37 ( .A(_647_), .B(_649_), .Y(_660_) );
	AOI22X1 AOI22X1_42 ( .A(_644_), .B(_660_), .C(_659_), .D(_640_), .Y(_661_) );
	NOR2X1 NOR2X1_231 ( .A(_642_), .B(_1068_), .Y(_662_) );
	OAI21X1 OAI21X1_398 ( .A(_633_), .B(_652_), .C(_662_), .Y(_663_) );
	INVX1 INVX1_136 ( .A(_663_), .Y(_664_) );
	NOR2X1 NOR2X1_232 ( .A(_885__bF_buf0), .B(_896__bF_buf0), .Y(_665_) );
	OAI22X1 OAI22X1_44 ( .A(_433_), .B(_1064_), .C(res), .D(_1057__bF_buf0), .Y(_666_) );
	AOI21X1 AOI21X1_95 ( .A(ABL_1_), .B(_665_), .C(_666_), .Y(_667_) );
	OAI21X1 OAI21X1_399 ( .A(_433_), .B(_627_), .C(_667_), .Y(_668_) );
	INVX1 INVX1_137 ( .A(_668_), .Y(_669_) );
	OAI21X1 OAI21X1_400 ( .A(_1418_), .B(_664_), .C(_669_), .Y(_670_) );
	NOR2X1 NOR2X1_233 ( .A(_661_), .B(_670_), .Y(_671_) );
	AOI21X1 AOI21X1_96 ( .A(_663_), .B(PC_1_), .C(_668_), .Y(_672_) );
	OAI21X1 OAI21X1_401 ( .A(_672_), .B(_657_), .C(RDY_bF_buf8), .Y(_673_) );
	OAI22X1 OAI22X1_45 ( .A(RDY_bF_buf7), .B(_1418_), .C(_673_), .D(_671_), .Y(_9__1_) );
	NOR2X1 NOR2X1_234 ( .A(_672_), .B(_657_), .Y(_674_) );
	AOI21X1 AOI21X1_97 ( .A(_632_), .B(_454_), .C(_115_), .Y(_675_) );
	NAND3X1 NAND3X1_112 ( .A(ADD_2_), .B(_882__bF_buf4), .C(_1034__bF_buf3), .Y(_676_) );
	NOR2X1 NOR2X1_235 ( .A(res), .B(_894_), .Y(_677_) );
	INVX1 INVX1_138 ( .A(_677_), .Y(_678_) );
	NAND3X1 NAND3X1_113 ( .A(_882__bF_buf3), .B(_678_), .C(_1046_), .Y(_679_) );
	NAND3X1 NAND3X1_114 ( .A(PC_2_), .B(_882__bF_buf2), .C(_483_), .Y(_680_) );
	NAND3X1 NAND3X1_115 ( .A(_680_), .B(_676_), .C(_679_), .Y(_681_) );
	NAND2X1 NAND2X1_191 ( .A(ABL_2_), .B(_910__bF_buf0), .Y(_682_) );
	OAI21X1 OAI21X1_402 ( .A(_1420_), .B(_910__bF_buf4), .C(_682_), .Y(_683_) );
	AND2X2 AND2X2_38 ( .A(_683_), .B(_1436_), .Y(_684_) );
	NOR3X1 NOR3X1_18 ( .A(_681_), .B(_675_), .C(_684_), .Y(_685_) );
	OAI21X1 OAI21X1_403 ( .A(_1420_), .B(_631_), .C(_685_), .Y(_686_) );
	NOR2X1 NOR2X1_236 ( .A(_686_), .B(_674_), .Y(_687_) );
	NOR3X1 NOR3X1_19 ( .A(_1420_), .B(_633_), .C(_652_), .Y(_688_) );
	OAI21X1 OAI21X1_404 ( .A(_625_), .B(_626_), .C(ADD_2_), .Y(_689_) );
	OAI22X1 OAI22X1_46 ( .A(_115_), .B(_1064_), .C(_1057__bF_buf3), .D(_677_), .Y(_690_) );
	AOI21X1 AOI21X1_98 ( .A(PC_2_), .B(_1068_), .C(_690_), .Y(_691_) );
	NAND2X1 NAND2X1_192 ( .A(_1436_), .B(_683_), .Y(_692_) );
	NAND3X1 NAND3X1_116 ( .A(_692_), .B(_691_), .C(_689_), .Y(_693_) );
	OAI21X1 OAI21X1_405 ( .A(_688_), .B(_693_), .C(_674_), .Y(_694_) );
	NAND2X1 NAND2X1_193 ( .A(RDY_bF_buf6), .B(_694_), .Y(_695_) );
	OAI22X1 OAI22X1_47 ( .A(RDY_bF_buf5), .B(_1420_), .C(_687_), .D(_695_), .Y(_9__2_) );
	AOI21X1 AOI21X1_99 ( .A(_632_), .B(_454_), .C(_199_), .Y(_696_) );
	NAND3X1 NAND3X1_117 ( .A(ADD_3_), .B(_882__bF_buf1), .C(_1034__bF_buf2), .Y(_697_) );
	NAND3X1 NAND3X1_118 ( .A(PC_3_), .B(_882__bF_buf0), .C(_483_), .Y(_698_) );
	NAND3X1 NAND3X1_119 ( .A(_1057__bF_buf2), .B(_698_), .C(_697_), .Y(_699_) );
	NAND2X1 NAND2X1_194 ( .A(PC_3_), .B(_896__bF_buf3), .Y(_700_) );
	NAND2X1 NAND2X1_195 ( .A(ABL_3_), .B(_910__bF_buf3), .Y(_701_) );
	AOI21X1 AOI21X1_100 ( .A(_700_), .B(_701_), .C(_885__bF_buf4), .Y(_702_) );
	NOR3X1 NOR3X1_20 ( .A(_702_), .B(_699_), .C(_696_), .Y(_703_) );
	OAI21X1 OAI21X1_406 ( .A(_1421_), .B(_631_), .C(_703_), .Y(_704_) );
	AOI21X1 AOI21X1_101 ( .A(_674_), .B(_686_), .C(_704_), .Y(_705_) );
	NAND3X1 NAND3X1_120 ( .A(PC_2_), .B(_627_), .C(_630_), .Y(_706_) );
	NAND3X1 NAND3X1_121 ( .A(PC_3_), .B(_627_), .C(_630_), .Y(_707_) );
	AOI22X1 AOI22X1_43 ( .A(_703_), .B(_707_), .C(_706_), .D(_685_), .Y(_708_) );
	NAND3X1 NAND3X1_122 ( .A(_708_), .B(_661_), .C(_670_), .Y(_709_) );
	NAND2X1 NAND2X1_196 ( .A(RDY_bF_buf4), .B(_709_), .Y(_710_) );
	OAI22X1 OAI22X1_48 ( .A(RDY_bF_buf3), .B(_1421_), .C(_710_), .D(_705_), .Y(_9__3_) );
	NOR3X1 NOR3X1_21 ( .A(_1421_), .B(_633_), .C(_652_), .Y(_711_) );
	OAI21X1 OAI21X1_407 ( .A(_625_), .B(_626_), .C(ADD_3_), .Y(_712_) );
	OAI21X1 OAI21X1_408 ( .A(_199_), .B(_1064_), .C(_1057__bF_buf1), .Y(_713_) );
	AOI21X1 AOI21X1_102 ( .A(PC_3_), .B(_1068_), .C(_713_), .Y(_714_) );
	OAI21X1 OAI21X1_409 ( .A(_1421_), .B(_910__bF_buf2), .C(_701_), .Y(_715_) );
	NAND2X1 NAND2X1_197 ( .A(_1436_), .B(_715_), .Y(_716_) );
	NAND3X1 NAND3X1_123 ( .A(_716_), .B(_714_), .C(_712_), .Y(_717_) );
	OAI22X1 OAI22X1_49 ( .A(_711_), .B(_717_), .C(_688_), .D(_693_), .Y(_718_) );
	NOR3X1 NOR3X1_22 ( .A(_672_), .B(_657_), .C(_718_), .Y(_719_) );
	AOI21X1 AOI21X1_103 ( .A(_632_), .B(_454_), .C(_551_), .Y(_720_) );
	NAND3X1 NAND3X1_124 ( .A(ADD_4_), .B(_882__bF_buf5), .C(_1034__bF_buf1), .Y(_721_) );
	NAND3X1 NAND3X1_125 ( .A(PC_4_), .B(_882__bF_buf4), .C(_483_), .Y(_722_) );
	NAND3X1 NAND3X1_126 ( .A(_1057__bF_buf0), .B(_722_), .C(_721_), .Y(_723_) );
	NAND2X1 NAND2X1_198 ( .A(PC_4_), .B(_896__bF_buf2), .Y(_724_) );
	NAND2X1 NAND2X1_199 ( .A(ABL_4_), .B(_910__bF_buf1), .Y(_725_) );
	AOI21X1 AOI21X1_104 ( .A(_724_), .B(_725_), .C(_885__bF_buf3), .Y(_726_) );
	NOR3X1 NOR3X1_23 ( .A(_726_), .B(_723_), .C(_720_), .Y(_727_) );
	OAI21X1 OAI21X1_410 ( .A(_1422_), .B(_631_), .C(_727_), .Y(_728_) );
	NOR2X1 NOR2X1_237 ( .A(_728_), .B(_719_), .Y(_729_) );
	INVX1 INVX1_139 ( .A(_728_), .Y(_730_) );
	OAI21X1 OAI21X1_411 ( .A(_730_), .B(_709_), .C(RDY_bF_buf2), .Y(_731_) );
	OAI22X1 OAI22X1_50 ( .A(RDY_bF_buf1), .B(_1422_), .C(_731_), .D(_729_), .Y(_9__4_) );
	AOI21X1 AOI21X1_105 ( .A(_632_), .B(_454_), .C(_209_), .Y(_732_) );
	NAND3X1 NAND3X1_127 ( .A(ADD_5_), .B(_882__bF_buf3), .C(_1034__bF_buf0), .Y(_733_) );
	NAND3X1 NAND3X1_128 ( .A(PC_5_), .B(_882__bF_buf2), .C(_483_), .Y(_734_) );
	NAND3X1 NAND3X1_129 ( .A(_1057__bF_buf3), .B(_734_), .C(_733_), .Y(_735_) );
	NAND2X1 NAND2X1_200 ( .A(PC_5_), .B(_896__bF_buf1), .Y(_736_) );
	NAND2X1 NAND2X1_201 ( .A(ABL_5_), .B(_910__bF_buf0), .Y(_737_) );
	AOI21X1 AOI21X1_106 ( .A(_736_), .B(_737_), .C(_885__bF_buf2), .Y(_738_) );
	NOR3X1 NOR3X1_24 ( .A(_738_), .B(_735_), .C(_732_), .Y(_739_) );
	OAI21X1 OAI21X1_412 ( .A(_1423_), .B(_631_), .C(_739_), .Y(_740_) );
	AOI21X1 AOI21X1_107 ( .A(_719_), .B(_728_), .C(_740_), .Y(_741_) );
	NAND3X1 NAND3X1_130 ( .A(PC_4_), .B(_627_), .C(_630_), .Y(_742_) );
	NAND3X1 NAND3X1_131 ( .A(PC_5_), .B(_627_), .C(_630_), .Y(_743_) );
	AOI22X1 AOI22X1_44 ( .A(_727_), .B(_742_), .C(_743_), .D(_739_), .Y(_744_) );
	INVX1 INVX1_140 ( .A(_744_), .Y(_745_) );
	OAI21X1 OAI21X1_413 ( .A(_745_), .B(_709_), .C(RDY_bF_buf0), .Y(_746_) );
	OAI22X1 OAI22X1_51 ( .A(RDY_bF_buf8), .B(_1423_), .C(_746_), .D(_741_), .Y(_9__5_) );
	AOI21X1 AOI21X1_108 ( .A(_632_), .B(_454_), .C(_224_), .Y(_747_) );
	NAND3X1 NAND3X1_132 ( .A(ADD_6_), .B(_882__bF_buf1), .C(_1034__bF_buf3), .Y(_748_) );
	NAND3X1 NAND3X1_133 ( .A(PC_6_), .B(_882__bF_buf0), .C(_483_), .Y(_749_) );
	NAND3X1 NAND3X1_134 ( .A(_1057__bF_buf2), .B(_749_), .C(_748_), .Y(_750_) );
	NAND2X1 NAND2X1_202 ( .A(PC_6_), .B(_896__bF_buf0), .Y(_751_) );
	NAND2X1 NAND2X1_203 ( .A(ABL_6_), .B(_910__bF_buf4), .Y(_752_) );
	AOI21X1 AOI21X1_109 ( .A(_751_), .B(_752_), .C(_885__bF_buf1), .Y(_753_) );
	NOR3X1 NOR3X1_25 ( .A(_753_), .B(_750_), .C(_747_), .Y(_754_) );
	OAI21X1 OAI21X1_414 ( .A(_1425_), .B(_631_), .C(_754_), .Y(_755_) );
	AOI21X1 AOI21X1_110 ( .A(_719_), .B(_744_), .C(_755_), .Y(_756_) );
	NAND3X1 NAND3X1_135 ( .A(_744_), .B(_755_), .C(_719_), .Y(_757_) );
	NAND2X1 NAND2X1_204 ( .A(RDY_bF_buf7), .B(_757_), .Y(_758_) );
	OAI22X1 OAI22X1_52 ( .A(RDY_bF_buf6), .B(_1425_), .C(_756_), .D(_758_), .Y(_9__6_) );
	AOI21X1 AOI21X1_111 ( .A(_632_), .B(_454_), .C(_421_), .Y(_759_) );
	NAND3X1 NAND3X1_136 ( .A(ADD_7_), .B(_882__bF_buf5), .C(_1034__bF_buf2), .Y(_760_) );
	NAND3X1 NAND3X1_137 ( .A(PC_7_), .B(_882__bF_buf4), .C(_483_), .Y(_761_) );
	NAND3X1 NAND3X1_138 ( .A(_1057__bF_buf1), .B(_761_), .C(_760_), .Y(_762_) );
	MUX2X1 MUX2X1_15 ( .A(ABL_7_), .B(PC_7_), .S(_910__bF_buf3), .Y(_763_) );
	NOR2X1 NOR2X1_238 ( .A(_885__bF_buf0), .B(_763_), .Y(_764_) );
	NOR3X1 NOR3X1_26 ( .A(_762_), .B(_764_), .C(_759_), .Y(_765_) );
	OAI21X1 OAI21X1_415 ( .A(_1426_), .B(_631_), .C(_765_), .Y(_766_) );
	INVX1 INVX1_141 ( .A(_766_), .Y(_767_) );
	AND2X2 AND2X2_39 ( .A(_757_), .B(_767_), .Y(_768_) );
	NAND3X1 NAND3X1_139 ( .A(PC_6_), .B(_627_), .C(_630_), .Y(_769_) );
	NAND3X1 NAND3X1_140 ( .A(PC_7_), .B(_627_), .C(_630_), .Y(_770_) );
	AOI22X1 AOI22X1_45 ( .A(_754_), .B(_769_), .C(_770_), .D(_765_), .Y(_771_) );
	NAND2X1 NAND2X1_205 ( .A(_744_), .B(_771_), .Y(_772_) );
	OAI21X1 OAI21X1_416 ( .A(_772_), .B(_709_), .C(RDY_bF_buf5), .Y(_773_) );
	OAI22X1 OAI22X1_53 ( .A(RDY_bF_buf4), .B(_1426_), .C(_773_), .D(_768_), .Y(_9__7_) );
	NAND2X1 NAND2X1_206 ( .A(PC_8_), .B(_881__bF_buf4), .Y(_774_) );
	NOR2X1 NOR2X1_239 ( .A(_772_), .B(_709_), .Y(_775_) );
	AOI21X1 AOI21X1_112 ( .A(_632_), .B(_454_), .C(_1403_), .Y(_776_) );
	NAND3X1 NAND3X1_141 ( .A(ADD_0_), .B(_882__bF_buf3), .C(_483_), .Y(_777_) );
	NAND3X1 NAND3X1_142 ( .A(_1057__bF_buf0), .B(_777_), .C(_1433_), .Y(_778_) );
	NAND2X1 NAND2X1_207 ( .A(PC_8_), .B(_896__bF_buf3), .Y(_779_) );
	NAND2X1 NAND2X1_208 ( .A(ABH_0_), .B(_910__bF_buf2), .Y(_780_) );
	AOI21X1 AOI21X1_113 ( .A(_779_), .B(_780_), .C(_885__bF_buf4), .Y(_781_) );
	NOR3X1 NOR3X1_27 ( .A(_781_), .B(_778_), .C(_776_), .Y(_782_) );
	OAI21X1 OAI21X1_417 ( .A(_102_), .B(_631_), .C(_782_), .Y(_783_) );
	XNOR2X1 XNOR2X1_8 ( .A(_775_), .B(_783_), .Y(_784_) );
	OAI21X1 OAI21X1_418 ( .A(_881__bF_buf3), .B(_784_), .C(_774_), .Y(_9__8_) );
	AOI21X1 AOI21X1_114 ( .A(_632_), .B(_454_), .C(_1419_), .Y(_785_) );
	NAND3X1 NAND3X1_143 ( .A(ADD_1_), .B(_882__bF_buf2), .C(_483_), .Y(_786_) );
	NAND3X1 NAND3X1_144 ( .A(_1057__bF_buf3), .B(_786_), .C(_1486_), .Y(_787_) );
	MUX2X1 MUX2X1_16 ( .A(ABH_1_), .B(PC_9_), .S(_910__bF_buf1), .Y(_788_) );
	NOR2X1 NOR2X1_240 ( .A(_885__bF_buf3), .B(_788_), .Y(_789_) );
	NOR3X1 NOR3X1_28 ( .A(_787_), .B(_789_), .C(_785_), .Y(_790_) );
	OAI21X1 OAI21X1_419 ( .A(_107_), .B(_631_), .C(_790_), .Y(_791_) );
	AOI21X1 AOI21X1_115 ( .A(_775_), .B(_783_), .C(_791_), .Y(_792_) );
	AND2X2 AND2X2_40 ( .A(_744_), .B(_771_), .Y(_793_) );
	NAND3X1 NAND3X1_145 ( .A(PC_8_), .B(_627_), .C(_630_), .Y(_794_) );
	NAND3X1 NAND3X1_146 ( .A(PC_9_), .B(_627_), .C(_630_), .Y(_795_) );
	AOI22X1 AOI22X1_46 ( .A(_782_), .B(_794_), .C(_795_), .D(_790_), .Y(_796_) );
	NAND3X1 NAND3X1_147 ( .A(_793_), .B(_796_), .C(_719_), .Y(_797_) );
	NAND2X1 NAND2X1_209 ( .A(RDY_bF_buf3), .B(_797_), .Y(_798_) );
	OAI22X1 OAI22X1_54 ( .A(RDY_bF_buf2), .B(_107_), .C(_798_), .D(_792_), .Y(_9__9_) );
	INVX1 INVX1_142 ( .A(_797_), .Y(_799_) );
	AOI21X1 AOI21X1_116 ( .A(_632_), .B(_454_), .C(_905_), .Y(_800_) );
	NAND3X1 NAND3X1_148 ( .A(ADD_2_), .B(_882__bF_buf1), .C(_483_), .Y(_801_) );
	NAND3X1 NAND3X1_149 ( .A(_1057__bF_buf2), .B(_801_), .C(_1498_), .Y(_802_) );
	NAND2X1 NAND2X1_210 ( .A(PC_10_), .B(_896__bF_buf2), .Y(_803_) );
	NAND2X1 NAND2X1_211 ( .A(ABH_2_), .B(_910__bF_buf0), .Y(_804_) );
	AOI21X1 AOI21X1_117 ( .A(_803_), .B(_804_), .C(_885__bF_buf2), .Y(_805_) );
	NOR3X1 NOR3X1_29 ( .A(_805_), .B(_802_), .C(_800_), .Y(_806_) );
	OAI21X1 OAI21X1_420 ( .A(_114_), .B(_631_), .C(_806_), .Y(_807_) );
	NOR2X1 NOR2X1_241 ( .A(_807_), .B(_799_), .Y(_808_) );
	INVX1 INVX1_143 ( .A(_807_), .Y(_809_) );
	OAI21X1 OAI21X1_421 ( .A(_809_), .B(_797_), .C(RDY_bF_buf1), .Y(_810_) );
	OAI22X1 OAI22X1_55 ( .A(RDY_bF_buf0), .B(_114_), .C(_810_), .D(_808_), .Y(_9__10_) );
	AOI21X1 AOI21X1_118 ( .A(_632_), .B(_454_), .C(_1095_), .Y(_811_) );
	NAND3X1 NAND3X1_150 ( .A(ADD_3_), .B(_882__bF_buf0), .C(_483_), .Y(_812_) );
	NAND3X1 NAND3X1_151 ( .A(_1057__bF_buf1), .B(_812_), .C(_1508_), .Y(_813_) );
	MUX2X1 MUX2X1_17 ( .A(ABH_3_), .B(PC_11_), .S(_910__bF_buf4), .Y(_814_) );
	NOR2X1 NOR2X1_242 ( .A(_885__bF_buf1), .B(_814_), .Y(_815_) );
	NOR3X1 NOR3X1_30 ( .A(_813_), .B(_815_), .C(_811_), .Y(_816_) );
	OAI21X1 OAI21X1_422 ( .A(_122_), .B(_631_), .C(_816_), .Y(_817_) );
	AOI21X1 AOI21X1_119 ( .A(_799_), .B(_807_), .C(_817_), .Y(_818_) );
	NAND3X1 NAND3X1_152 ( .A(PC_10_), .B(_627_), .C(_630_), .Y(_819_) );
	NAND3X1 NAND3X1_153 ( .A(PC_11_), .B(_627_), .C(_630_), .Y(_820_) );
	AOI22X1 AOI22X1_47 ( .A(_806_), .B(_819_), .C(_820_), .D(_816_), .Y(_821_) );
	INVX1 INVX1_144 ( .A(_821_), .Y(_822_) );
	OAI21X1 OAI21X1_423 ( .A(_822_), .B(_797_), .C(RDY_bF_buf8), .Y(_823_) );
	OAI22X1 OAI22X1_56 ( .A(RDY_bF_buf7), .B(_122_), .C(_823_), .D(_818_), .Y(_9__11_) );
	NOR2X1 NOR2X1_243 ( .A(_822_), .B(_797_), .Y(_824_) );
	NOR2X1 NOR2X1_244 ( .A(_131_), .B(_631_), .Y(_825_) );
	OAI21X1 OAI21X1_424 ( .A(_1525_), .B(_1064_), .C(_1057__bF_buf0), .Y(_826_) );
	AOI21X1 AOI21X1_120 ( .A(ADD_4_), .B(_1068_), .C(_826_), .Y(_827_) );
	NOR2X1 NOR2X1_245 ( .A(_131_), .B(_910__bF_buf3), .Y(_828_) );
	NOR2X1 NOR2X1_246 ( .A(_1525_), .B(_896__bF_buf1), .Y(_829_) );
	OAI21X1 OAI21X1_425 ( .A(_828_), .B(_829_), .C(_1436_), .Y(_830_) );
	AND2X2 AND2X2_41 ( .A(_827_), .B(_830_), .Y(_831_) );
	OAI21X1 OAI21X1_426 ( .A(_891_), .B(_627_), .C(_831_), .Y(_832_) );
	OR2X2 OR2X2_31 ( .A(_832_), .B(_825_), .Y(_833_) );
	NOR2X1 NOR2X1_247 ( .A(_833_), .B(_824_), .Y(_834_) );
	NAND3X1 NAND3X1_154 ( .A(_796_), .B(_821_), .C(_775_), .Y(_835_) );
	INVX1 INVX1_145 ( .A(_833_), .Y(_836_) );
	OAI21X1 OAI21X1_427 ( .A(_836_), .B(_835_), .C(RDY_bF_buf6), .Y(_837_) );
	OAI22X1 OAI22X1_57 ( .A(RDY_bF_buf5), .B(_131_), .C(_837_), .D(_834_), .Y(_9__12_) );
	NOR2X1 NOR2X1_248 ( .A(_633_), .B(_652_), .Y(_838_) );
	OAI21X1 OAI21X1_428 ( .A(_642_), .B(_838_), .C(PC_13_), .Y(_839_) );
	OAI21X1 OAI21X1_429 ( .A(_625_), .B(_626_), .C(DIMUX_5_), .Y(_840_) );
	INVX1 INVX1_146 ( .A(_1068_), .Y(_841_) );
	AOI21X1 AOI21X1_121 ( .A(_1224_), .B(ABH_5_), .C(_1194_), .Y(_842_) );
	OAI21X1 OAI21X1_430 ( .A(_209_), .B(_841_), .C(_842_), .Y(_843_) );
	AOI21X1 AOI21X1_122 ( .A(ABH_5_), .B(_665_), .C(_843_), .Y(_844_) );
	NAND3X1 NAND3X1_155 ( .A(_840_), .B(_844_), .C(_839_), .Y(_845_) );
	AOI21X1 AOI21X1_123 ( .A(_824_), .B(_833_), .C(_845_), .Y(_846_) );
	OAI21X1 OAI21X1_431 ( .A(_825_), .B(_832_), .C(_845_), .Y(_847_) );
	OAI21X1 OAI21X1_432 ( .A(_847_), .B(_835_), .C(RDY_bF_buf4), .Y(_848_) );
	OAI22X1 OAI22X1_58 ( .A(RDY_bF_buf3), .B(_135_), .C(_848_), .D(_846_), .Y(_9__13_) );
	NAND2X1 NAND2X1_212 ( .A(_796_), .B(_821_), .Y(_849_) );
	NOR3X1 NOR3X1_31 ( .A(_772_), .B(_849_), .C(_709_), .Y(_850_) );
	INVX1 INVX1_147 ( .A(_847_), .Y(_851_) );
	OAI21X1 OAI21X1_433 ( .A(_642_), .B(_838_), .C(PC_14_), .Y(_852_) );
	INVX1 INVX1_148 ( .A(_665_), .Y(_853_) );
	OAI21X1 OAI21X1_434 ( .A(_52_), .B(_1064_), .C(_1057__bF_buf3), .Y(_854_) );
	AOI21X1 AOI21X1_124 ( .A(ADD_6_), .B(_1068_), .C(_854_), .Y(_855_) );
	OAI21X1 OAI21X1_435 ( .A(_52_), .B(_853_), .C(_855_), .Y(_856_) );
	AOI21X1 AOI21X1_125 ( .A(DIMUX_6_), .B(_633_), .C(_856_), .Y(_857_) );
	AOI22X1 AOI22X1_48 ( .A(_852_), .B(_857_), .C(_851_), .D(_850_), .Y(_858_) );
	AND2X2 AND2X2_42 ( .A(_796_), .B(_821_), .Y(_859_) );
	NAND3X1 NAND3X1_156 ( .A(_793_), .B(_859_), .C(_719_), .Y(_860_) );
	NAND2X1 NAND2X1_213 ( .A(_852_), .B(_857_), .Y(_861_) );
	NOR3X1 NOR3X1_32 ( .A(_847_), .B(_861_), .C(_860_), .Y(_862_) );
	OAI21X1 OAI21X1_436 ( .A(_858_), .B(_862_), .C(RDY_bF_buf2), .Y(_863_) );
	OAI21X1 OAI21X1_437 ( .A(RDY_bF_buf1), .B(_142_), .C(_863_), .Y(_9__14_) );
	NOR3X1 NOR3X1_33 ( .A(_822_), .B(_847_), .C(_797_), .Y(_864_) );
	NOR2X1 NOR2X1_249 ( .A(_62_), .B(_853_), .Y(_865_) );
	OAI21X1 OAI21X1_438 ( .A(_642_), .B(_838_), .C(PC_15_), .Y(_866_) );
	OAI21X1 OAI21X1_439 ( .A(_625_), .B(_626_), .C(DIMUX_7_), .Y(_867_) );
	OAI21X1 OAI21X1_440 ( .A(_62_), .B(_1064_), .C(_1057__bF_buf2), .Y(_868_) );
	AOI21X1 AOI21X1_126 ( .A(ADD_7_), .B(_1068_), .C(_868_), .Y(_869_) );
	NAND3X1 NAND3X1_157 ( .A(_867_), .B(_869_), .C(_866_), .Y(_870_) );
	NOR2X1 NOR2X1_250 ( .A(_865_), .B(_870_), .Y(_871_) );
	NAND3X1 NAND3X1_158 ( .A(_861_), .B(_871_), .C(_864_), .Y(_872_) );
	INVX1 INVX1_149 ( .A(_871_), .Y(_873_) );
	NAND3X1 NAND3X1_159 ( .A(_851_), .B(_861_), .C(_850_), .Y(_874_) );
	AOI21X1 AOI21X1_127 ( .A(_874_), .B(_873_), .C(_881__bF_buf2), .Y(_875_) );
	AOI22X1 AOI22X1_49 ( .A(_881__bF_buf1), .B(_147_), .C(_872_), .D(_875_), .Y(_9__15_) );
	BUFX2 BUFX2_9 ( .A(_1536__0_), .Y(AB[0]) );
	BUFX2 BUFX2_10 ( .A(_1536__1_), .Y(AB[1]) );
	BUFX2 BUFX2_11 ( .A(_1536__2_), .Y(AB[2]) );
	BUFX2 BUFX2_12 ( .A(_1536__3_), .Y(AB[3]) );
	BUFX2 BUFX2_13 ( .A(_1536__4_), .Y(AB[4]) );
	BUFX2 BUFX2_14 ( .A(_1536__5_), .Y(AB[5]) );
	BUFX2 BUFX2_15 ( .A(_1536__6_), .Y(AB[6]) );
	BUFX2 BUFX2_16 ( .A(_1536__7_), .Y(AB[7]) );
	BUFX2 BUFX2_17 ( .A(_1536__8_), .Y(AB[8]) );
	BUFX2 BUFX2_18 ( .A(_1536__9_), .Y(AB[9]) );
	BUFX2 BUFX2_19 ( .A(_1536__10_), .Y(AB[10]) );
	BUFX2 BUFX2_20 ( .A(_1536__11_), .Y(AB[11]) );
	BUFX2 BUFX2_21 ( .A(_1536__12_), .Y(AB[12]) );
	BUFX2 BUFX2_22 ( .A(_1536__13_), .Y(AB[13]) );
	BUFX2 BUFX2_23 ( .A(_1536__14_), .Y(AB[14]) );
	BUFX2 BUFX2_24 ( .A(_1536__15_), .Y(AB[15]) );
	BUFX2 BUFX2_25 ( .A(_1537__0_), .Y(DO[0]) );
	BUFX2 BUFX2_26 ( .A(_1537__1_), .Y(DO[1]) );
	BUFX2 BUFX2_27 ( .A(_1537__2_), .Y(DO[2]) );
	BUFX2 BUFX2_28 ( .A(_1537__3_), .Y(DO[3]) );
	BUFX2 BUFX2_29 ( .A(_1537__4_), .Y(DO[4]) );
	BUFX2 BUFX2_30 ( .A(_1537__5_), .Y(DO[5]) );
	BUFX2 BUFX2_31 ( .A(_1537__6_), .Y(DO[6]) );
	BUFX2 BUFX2_32 ( .A(_1537__7_), .Y(DO[7]) );
	BUFX2 BUFX2_33 ( .A(_1538_), .Y(WE) );
	DFFPOSX1 DFFPOSX1_1 ( .CLK(clk_bF_buf11), .D(_1328_), .Q(AXYS_0__0_) );
	DFFPOSX1 DFFPOSX1_2 ( .CLK(clk_bF_buf10), .D(_1345_), .Q(AXYS_0__1_) );
	DFFPOSX1 DFFPOSX1_3 ( .CLK(clk_bF_buf9), .D(_1352_), .Q(AXYS_0__2_) );
	DFFPOSX1 DFFPOSX1_4 ( .CLK(clk_bF_buf8), .D(_1359_), .Q(AXYS_0__3_) );
	DFFPOSX1 DFFPOSX1_5 ( .CLK(clk_bF_buf7), .D(_1363_), .Q(AXYS_0__4_) );
	DFFPOSX1 DFFPOSX1_6 ( .CLK(clk_bF_buf6), .D(_1375_), .Q(AXYS_0__5_) );
	DFFPOSX1 DFFPOSX1_7 ( .CLK(clk_bF_buf5), .D(_1381_), .Q(AXYS_0__6_) );
	DFFPOSX1 DFFPOSX1_8 ( .CLK(clk_bF_buf4), .D(_1389_), .Q(AXYS_0__7_) );
	DFFPOSX1 DFFPOSX1_9 ( .CLK(clk_bF_buf3), .D(_68_), .Q(AXYS_1__0_) );
	DFFPOSX1 DFFPOSX1_10 ( .CLK(clk_bF_buf2), .D(_71_), .Q(AXYS_1__1_) );
	DFFPOSX1 DFFPOSX1_11 ( .CLK(clk_bF_buf1), .D(_74_), .Q(AXYS_1__2_) );
	DFFPOSX1 DFFPOSX1_12 ( .CLK(clk_bF_buf0), .D(_76_), .Q(AXYS_1__3_) );
	DFFPOSX1 DFFPOSX1_13 ( .CLK(clk_bF_buf11), .D(_79_), .Q(AXYS_1__4_) );
	DFFPOSX1 DFFPOSX1_14 ( .CLK(clk_bF_buf10), .D(_82_), .Q(AXYS_1__5_) );
	DFFPOSX1 DFFPOSX1_15 ( .CLK(clk_bF_buf9), .D(_84_), .Q(AXYS_1__6_) );
	DFFPOSX1 DFFPOSX1_16 ( .CLK(clk_bF_buf8), .D(_86_), .Q(AXYS_1__7_) );
	DFFPOSX1 DFFPOSX1_17 ( .CLK(clk_bF_buf7), .D(_153_), .Q(AXYS_3__0_) );
	DFFPOSX1 DFFPOSX1_18 ( .CLK(clk_bF_buf6), .D(_154_), .Q(AXYS_3__1_) );
	DFFPOSX1 DFFPOSX1_19 ( .CLK(clk_bF_buf5), .D(_156_), .Q(AXYS_3__2_) );
	DFFPOSX1 DFFPOSX1_20 ( .CLK(clk_bF_buf4), .D(_159_), .Q(AXYS_3__3_) );
	DFFPOSX1 DFFPOSX1_21 ( .CLK(clk_bF_buf3), .D(_162_), .Q(AXYS_3__4_) );
	DFFPOSX1 DFFPOSX1_22 ( .CLK(clk_bF_buf2), .D(_165_), .Q(AXYS_3__5_) );
	DFFPOSX1 DFFPOSX1_23 ( .CLK(clk_bF_buf1), .D(_168_), .Q(AXYS_3__6_) );
	DFFPOSX1 DFFPOSX1_24 ( .CLK(clk_bF_buf0), .D(_171_), .Q(AXYS_3__7_) );
	DFFPOSX1 DFFPOSX1_25 ( .CLK(clk_bF_buf11), .D(_1510_), .Q(AXYS_2__0_) );
	DFFPOSX1 DFFPOSX1_26 ( .CLK(clk_bF_buf10), .D(_1513_), .Q(AXYS_2__1_) );
	DFFPOSX1 DFFPOSX1_27 ( .CLK(clk_bF_buf9), .D(_1516_), .Q(AXYS_2__2_) );
	DFFPOSX1 DFFPOSX1_28 ( .CLK(clk_bF_buf8), .D(_1519_), .Q(AXYS_2__3_) );
	DFFPOSX1 DFFPOSX1_29 ( .CLK(clk_bF_buf7), .D(_1522_), .Q(AXYS_2__4_) );
	DFFPOSX1 DFFPOSX1_30 ( .CLK(clk_bF_buf6), .D(_1524_), .Q(AXYS_2__5_) );
	DFFPOSX1 DFFPOSX1_31 ( .CLK(clk_bF_buf5), .D(_1527_), .Q(AXYS_2__6_) );
	DFFPOSX1 DFFPOSX1_32 ( .CLK(clk_bF_buf4), .D(_1530_), .Q(AXYS_2__7_) );
	DFFPOSX1 DFFPOSX1_33 ( .CLK(clk_bF_buf3), .D(_7_), .Q(NMI_edge) );
	DFFPOSX1 DFFPOSX1_34 ( .CLK(clk_bF_buf2), .D(NMI), .Q(NMI_1) );
	DFFPOSX1 DFFPOSX1_35 ( .CLK(clk_bF_buf1), .D(_22__0_), .Q(cond_code_0_) );
	DFFPOSX1 DFFPOSX1_36 ( .CLK(clk_bF_buf0), .D(_22__1_), .Q(cond_code_1_) );
	DFFPOSX1 DFFPOSX1_37 ( .CLK(clk_bF_buf11), .D(_22__2_), .Q(cond_code_2_) );
	DFFPOSX1 DFFPOSX1_38 ( .CLK(clk_bF_buf10), .D(_30_), .Q(plp) );
	DFFPOSX1 DFFPOSX1_39 ( .CLK(clk_bF_buf9), .D(_29_), .Q(php) );
	DFFPOSX1 DFFPOSX1_40 ( .CLK(clk_bF_buf8), .D(_17_), .Q(clc) );
	DFFPOSX1 DFFPOSX1_41 ( .CLK(clk_bF_buf7), .D(_33_), .Q(sec) );
	DFFPOSX1 DFFPOSX1_42 ( .CLK(clk_bF_buf6), .D(_18_), .Q(cld) );
	DFFPOSX1 DFFPOSX1_43 ( .CLK(clk_bF_buf5), .D(_34_), .Q(sed) );
	DFFPOSX1 DFFPOSX1_44 ( .CLK(clk_bF_buf4), .D(_19_), .Q(cli) );
	DFFPOSX1 DFFPOSX1_45 ( .CLK(clk_bF_buf3), .D(_35_), .Q(sei) );
	DFFPOSX1 DFFPOSX1_46 ( .CLK(clk_bF_buf2), .D(_20_), .Q(clv) );
	DFFPOSX1 DFFPOSX1_47 ( .CLK(clk_bF_buf1), .D(_16_), .Q(bit_ins) );
	DFFPOSX1 DFFPOSX1_48 ( .CLK(clk_bF_buf0), .D(_28__0_), .Q(op_0_) );
	DFFPOSX1 DFFPOSX1_49 ( .CLK(clk_bF_buf11), .D(_28__1_), .Q(op_1_) );
	DFFPOSX1 DFFPOSX1_50 ( .CLK(clk_bF_buf10), .D(_28__2_), .Q(op_2_) );
	DFFPOSX1 DFFPOSX1_51 ( .CLK(clk_bF_buf9), .D(_28__3_), .Q(op_3_) );
	DFFPOSX1 DFFPOSX1_52 ( .CLK(clk_bF_buf8), .D(_32_), .Q(rotate) );
	DFFPOSX1 DFFPOSX1_53 ( .CLK(clk_bF_buf7), .D(_37_), .Q(shift_right) );
	DFFPOSX1 DFFPOSX1_54 ( .CLK(clk_bF_buf6), .D(_21_), .Q(compare) );
	DFFPOSX1 DFFPOSX1_55 ( .CLK(clk_bF_buf5), .D(_36_), .Q(shift) );
	DFFPOSX1 DFFPOSX1_56 ( .CLK(clk_bF_buf4), .D(_12_), .Q(adc_bcd) );
	DFFPOSX1 DFFPOSX1_57 ( .CLK(clk_bF_buf3), .D(_13_), .Q(adc_sbc) );
	DFFPOSX1 DFFPOSX1_58 ( .CLK(clk_bF_buf2), .D(_24_), .Q(inc) );
	DFFPOSX1 DFFPOSX1_59 ( .CLK(clk_bF_buf1), .D(_26_), .Q(load_only) );
	DFFPOSX1 DFFPOSX1_60 ( .CLK(clk_bF_buf0), .D(_40_), .Q(write_back) );
	DFFPOSX1 DFFPOSX1_61 ( .CLK(clk_bF_buf11), .D(_39_), .Q(store) );
	DFFPOSX1 DFFPOSX1_62 ( .CLK(clk_bF_buf10), .D(_25_), .Q(index_y) );
	DFFPOSX1 DFFPOSX1_63 ( .CLK(clk_bF_buf9), .D(_38__0_), .Q(src_reg_0_) );
	DFFPOSX1 DFFPOSX1_64 ( .CLK(clk_bF_buf8), .D(_38__1_), .Q(src_reg_1_) );
	DFFPOSX1 DFFPOSX1_65 ( .CLK(clk_bF_buf7), .D(_23__0_), .Q(dst_reg_0_) );
	DFFPOSX1 DFFPOSX1_66 ( .CLK(clk_bF_buf6), .D(_23__1_), .Q(dst_reg_1_) );
	DFFPOSX1 DFFPOSX1_67 ( .CLK(clk_bF_buf5), .D(_27_), .Q(load_reg) );
	DFFPOSX1 DFFPOSX1_68 ( .CLK(clk_bF_buf4), .D(_31_), .Q(res) );
	DFFPOSX1 DFFPOSX1_69 ( .CLK(clk_bF_buf3), .D(DIMUX_0_), .Q(DIHOLD_0_) );
	DFFPOSX1 DFFPOSX1_70 ( .CLK(clk_bF_buf2), .D(DIMUX_1_), .Q(DIHOLD_1_) );
	DFFPOSX1 DFFPOSX1_71 ( .CLK(clk_bF_buf1), .D(DIMUX_2_), .Q(DIHOLD_2_) );
	DFFPOSX1 DFFPOSX1_72 ( .CLK(clk_bF_buf0), .D(DIMUX_3_), .Q(DIHOLD_3_) );
	DFFPOSX1 DFFPOSX1_73 ( .CLK(clk_bF_buf11), .D(DIMUX_4_), .Q(DIHOLD_4_) );
	DFFPOSX1 DFFPOSX1_74 ( .CLK(clk_bF_buf10), .D(DIMUX_5_), .Q(DIHOLD_5_) );
	DFFPOSX1 DFFPOSX1_75 ( .CLK(clk_bF_buf9), .D(DIMUX_6_), .Q(DIHOLD_6_) );
	DFFPOSX1 DFFPOSX1_76 ( .CLK(clk_bF_buf8), .D(DIMUX_7_), .Q(DIHOLD_7_) );
	DFFPOSX1 DFFPOSX1_77 ( .CLK(clk_bF_buf7), .D(_4__0_), .Q(IRHOLD_0_) );
	DFFPOSX1 DFFPOSX1_78 ( .CLK(clk_bF_buf6), .D(_4__1_), .Q(IRHOLD_1_) );
	DFFPOSX1 DFFPOSX1_79 ( .CLK(clk_bF_buf5), .D(_4__2_), .Q(IRHOLD_2_) );
	DFFPOSX1 DFFPOSX1_80 ( .CLK(clk_bF_buf4), .D(_4__3_), .Q(IRHOLD_3_) );
	DFFPOSX1 DFFPOSX1_81 ( .CLK(clk_bF_buf3), .D(_4__4_), .Q(IRHOLD_4_) );
	DFFPOSX1 DFFPOSX1_82 ( .CLK(clk_bF_buf2), .D(_4__5_), .Q(IRHOLD_5_) );
	DFFPOSX1 DFFPOSX1_83 ( .CLK(clk_bF_buf1), .D(_4__6_), .Q(IRHOLD_6_) );
	DFFPOSX1 DFFPOSX1_84 ( .CLK(clk_bF_buf0), .D(_4__7_), .Q(IRHOLD_7_) );
	DFFPOSX1 DFFPOSX1_85 ( .CLK(clk_bF_buf11), .D(_5_), .Q(IRHOLD_valid) );
	DFFPOSX1 DFFPOSX1_86 ( .CLK(clk_bF_buf10), .D(_10_), .Q(V) );
	DFFPOSX1 DFFPOSX1_87 ( .CLK(clk_bF_buf9), .D(_3_), .Q(D) );
	DFFPOSX1 DFFPOSX1_88 ( .CLK(clk_bF_buf8), .D(_6_), .Q(I) );
	DFFPOSX1 DFFPOSX1_89 ( .CLK(clk_bF_buf7), .D(_8_), .Q(N) );
	DFFPOSX1 DFFPOSX1_90 ( .CLK(clk_bF_buf6), .D(_11_), .Q(Z) );
	DFFPOSX1 DFFPOSX1_91 ( .CLK(clk_bF_buf5), .D(_2_), .Q(C) );
	DFFPOSX1 DFFPOSX1_92 ( .CLK(clk_bF_buf4), .D(_15_), .Q(backwards) );
	DFFPOSX1 DFFPOSX1_93 ( .CLK(clk_bF_buf3), .D(_14_), .Q(adj_bcd) );
	DFFPOSX1 DFFPOSX1_94 ( .CLK(clk_bF_buf2), .D(_1__0_), .Q(ABL_0_) );
	DFFPOSX1 DFFPOSX1_95 ( .CLK(clk_bF_buf1), .D(_1__1_), .Q(ABL_1_) );
	DFFPOSX1 DFFPOSX1_96 ( .CLK(clk_bF_buf0), .D(_1__2_), .Q(ABL_2_) );
	DFFPOSX1 DFFPOSX1_97 ( .CLK(clk_bF_buf11), .D(_1__3_), .Q(ABL_3_) );
	DFFPOSX1 DFFPOSX1_98 ( .CLK(clk_bF_buf10), .D(_1__4_), .Q(ABL_4_) );
	DFFPOSX1 DFFPOSX1_99 ( .CLK(clk_bF_buf9), .D(_1__5_), .Q(ABL_5_) );
	DFFPOSX1 DFFPOSX1_100 ( .CLK(clk_bF_buf8), .D(_1__6_), .Q(ABL_6_) );
	DFFPOSX1 DFFPOSX1_101 ( .CLK(clk_bF_buf7), .D(_1__7_), .Q(ABL_7_) );
	DFFPOSX1 DFFPOSX1_102 ( .CLK(clk_bF_buf6), .D(_0__0_), .Q(ABH_0_) );
	DFFPOSX1 DFFPOSX1_103 ( .CLK(clk_bF_buf5), .D(_0__1_), .Q(ABH_1_) );
	DFFPOSX1 DFFPOSX1_104 ( .CLK(clk_bF_buf4), .D(_0__2_), .Q(ABH_2_) );
	DFFPOSX1 DFFPOSX1_105 ( .CLK(clk_bF_buf3), .D(_0__3_), .Q(ABH_3_) );
	DFFPOSX1 DFFPOSX1_106 ( .CLK(clk_bF_buf2), .D(_0__4_), .Q(ABH_4_) );
	DFFPOSX1 DFFPOSX1_107 ( .CLK(clk_bF_buf1), .D(_0__5_), .Q(ABH_5_) );
	DFFPOSX1 DFFPOSX1_108 ( .CLK(clk_bF_buf0), .D(_0__6_), .Q(ABH_6_) );
	DFFPOSX1 DFFPOSX1_109 ( .CLK(clk_bF_buf11), .D(_0__7_), .Q(ABH_7_) );
	DFFPOSX1 DFFPOSX1_110 ( .CLK(clk_bF_buf10), .D(_9__0_), .Q(PC_0_) );
	DFFPOSX1 DFFPOSX1_111 ( .CLK(clk_bF_buf9), .D(_9__1_), .Q(PC_1_) );
	DFFPOSX1 DFFPOSX1_112 ( .CLK(clk_bF_buf8), .D(_9__2_), .Q(PC_2_) );
	DFFPOSX1 DFFPOSX1_113 ( .CLK(clk_bF_buf7), .D(_9__3_), .Q(PC_3_) );
	DFFPOSX1 DFFPOSX1_114 ( .CLK(clk_bF_buf6), .D(_9__4_), .Q(PC_4_) );
	DFFPOSX1 DFFPOSX1_115 ( .CLK(clk_bF_buf5), .D(_9__5_), .Q(PC_5_) );
	DFFPOSX1 DFFPOSX1_116 ( .CLK(clk_bF_buf4), .D(_9__6_), .Q(PC_6_) );
	DFFPOSX1 DFFPOSX1_117 ( .CLK(clk_bF_buf3), .D(_9__7_), .Q(PC_7_) );
	DFFPOSX1 DFFPOSX1_118 ( .CLK(clk_bF_buf2), .D(_9__8_), .Q(PC_8_) );
	DFFPOSX1 DFFPOSX1_119 ( .CLK(clk_bF_buf1), .D(_9__9_), .Q(PC_9_) );
	DFFPOSX1 DFFPOSX1_120 ( .CLK(clk_bF_buf0), .D(_9__10_), .Q(PC_10_) );
	DFFPOSX1 DFFPOSX1_121 ( .CLK(clk_bF_buf11), .D(_9__11_), .Q(PC_11_) );
	DFFPOSX1 DFFPOSX1_122 ( .CLK(clk_bF_buf10), .D(_9__12_), .Q(PC_12_) );
	DFFPOSX1 DFFPOSX1_123 ( .CLK(clk_bF_buf9), .D(_9__13_), .Q(PC_13_) );
	DFFPOSX1 DFFPOSX1_124 ( .CLK(clk_bF_buf8), .D(_9__14_), .Q(PC_14_) );
	DFFPOSX1 DFFPOSX1_125 ( .CLK(clk_bF_buf7), .D(_9__15_), .Q(PC_15_) );
	DFFSR DFFSR_1 ( .CLK(clk_bF_buf6), .D(_876_), .Q(state_0_), .R(_1214_), .S(vdd) );
	DFFSR DFFSR_2 ( .CLK(clk_bF_buf5), .D(_877_), .Q(state_1_), .R(_1214_), .S(vdd) );
	DFFSR DFFSR_3 ( .CLK(clk_bF_buf4), .D(_878_), .Q(state_2_), .R(_1214_), .S(vdd) );
	DFFSR DFFSR_4 ( .CLK(clk_bF_buf3), .D(_879_), .Q(state_3_), .R(vdd), .S(_1214_) );
	DFFSR DFFSR_5 ( .CLK(clk_bF_buf2), .D(_880_), .Q(state_4_), .R(_1214_), .S(vdd) );
	DFFSR DFFSR_6 ( .CLK(clk_bF_buf1), .D(_888_), .Q(state_5_), .R(_1214_), .S(vdd) );
	OR2X2 OR2X2_32 ( .A(ADD_3_), .B(ADD_0_), .Y(_1711_) );
	NOR2X1 NOR2X1_251 ( .A(ADD_6_), .B(ADD_7_), .Y(_1712_) );
	NOR2X1 NOR2X1_252 ( .A(ADD_4_), .B(ADD_5_), .Y(_1713_) );
	NOR2X1 NOR2X1_253 ( .A(ADD_2_), .B(ADD_1_), .Y(_1714_) );
	NAND3X1 NAND3X1_160 ( .A(_1712_), .B(_1713_), .C(_1714_), .Y(_1715_) );
	NOR2X1 NOR2X1_254 ( .A(_1711_), .B(_1715_), .Y(ALU_Z) );
	INVX1 INVX1_150 ( .A(AI_7_), .Y(_1716_) );
	INVX8 INVX8_6 ( .A(RDY_bF_buf0), .Y(_1717_) );
	NAND2X1 NAND2X1_214 ( .A(ALU_AI7), .B(_1717__bF_buf3), .Y(_1718_) );
	OAI21X1 OAI21X1_441 ( .A(_1716_), .B(_1717__bF_buf2), .C(_1718_), .Y(_1539_) );
	NAND2X1 NAND2X1_215 ( .A(ALU_CI), .B(ALU_right), .Y(_1719_) );
	INVX4 INVX4_16 ( .A(ALU_op_1_), .Y(_1720_) );
	NAND2X1 NAND2X1_216 ( .A(ALU_op_0_), .B(_1720_), .Y(_1721_) );
	INVX2 INVX2_39 ( .A(ALU_op_0_), .Y(_1722_) );
	AND2X2 AND2X2_43 ( .A(_1722_), .B(ALU_BI_7_), .Y(_1723_) );
	NAND2X1 NAND2X1_217 ( .A(AI_7_), .B(_1723_), .Y(_1724_) );
	AOI22X1 AOI22X1_50 ( .A(ALU_BI_7_), .B(_1720_), .C(_1721_), .D(_1724_), .Y(_1725_) );
	INVX4 INVX4_17 ( .A(ALU_right), .Y(_1726_) );
	OAI21X1 OAI21X1_442 ( .A(AI_7_), .B(_1723_), .C(_1726_), .Y(_1727_) );
	OAI21X1 OAI21X1_443 ( .A(_1727_), .B(_1725_), .C(_1719_), .Y(_1728_) );
	INVX2 INVX2_40 ( .A(ALU_op_2_), .Y(_1729_) );
	NOR2X1 NOR2X1_255 ( .A(ALU_op_3_), .B(_1729_), .Y(_1730_) );
	INVX2 INVX2_41 ( .A(_1730_), .Y(_1731_) );
	NOR2X1 NOR2X1_256 ( .A(ALU_BI_7_), .B(_1731_), .Y(_1732_) );
	NOR2X1 NOR2X1_257 ( .A(ALU_op_3_), .B(ALU_op_2_), .Y(_1733_) );
	AOI21X1 AOI21X1_128 ( .A(ALU_BI_7_), .B(_1733_), .C(_1732_), .Y(_1734_) );
	INVX1 INVX1_151 ( .A(_1734_), .Y(_1735_) );
	INVX4 INVX4_18 ( .A(ALU_op_3_), .Y(_1736_) );
	OAI21X1 OAI21X1_444 ( .A(_1736_), .B(ALU_op_2_), .C(_1734_), .Y(_1737_) );
	OAI21X1 OAI21X1_445 ( .A(_1728_), .B(_1735_), .C(_1737_), .Y(_1738_) );
	NAND2X1 NAND2X1_218 ( .A(ALU_BI7), .B(_1717__bF_buf1), .Y(_1739_) );
	OAI21X1 OAI21X1_446 ( .A(_1717__bF_buf0), .B(_1738_), .C(_1739_), .Y(_1540_) );
	NAND2X1 NAND2X1_219 ( .A(ADD_0_), .B(_1717__bF_buf3), .Y(_1740_) );
	OAI21X1 OAI21X1_447 ( .A(_1736_), .B(_1729_), .C(ALU_CI), .Y(_1741_) );
	NOR2X1 NOR2X1_258 ( .A(ALU_right), .B(_1741_), .Y(_1742_) );
	NOR2X1 NOR2X1_259 ( .A(ALU_op_2_), .B(_1736_), .Y(_1743_) );
	NAND2X1 NAND2X1_220 ( .A(ALU_BI_0_), .B(_1722_), .Y(_1744_) );
	NAND2X1 NAND2X1_221 ( .A(ALU_op_1_), .B(AI_0_), .Y(_1745_) );
	AOI22X1 AOI22X1_51 ( .A(ALU_BI_0_), .B(_1745_), .C(_1721_), .D(_1744_), .Y(_1746_) );
	INVX1 INVX1_152 ( .A(ALU_BI_0_), .Y(_1747_) );
	INVX1 INVX1_153 ( .A(AI_0_), .Y(_1748_) );
	OAI21X1 OAI21X1_448 ( .A(ALU_op_0_), .B(_1747_), .C(_1748_), .Y(_1749_) );
	NAND2X1 NAND2X1_222 ( .A(_1726_), .B(_1749_), .Y(_1750_) );
	NAND2X1 NAND2X1_223 ( .A(ALU_right), .B(AI_1_), .Y(_1751_) );
	OAI21X1 OAI21X1_449 ( .A(_1746_), .B(_1750_), .C(_1751_), .Y(_1752_) );
	MUX2X1 MUX2X1_18 ( .A(_1730_), .B(_1733_), .S(_1747_), .Y(_1753_) );
	INVX1 INVX1_154 ( .A(_1753_), .Y(_1754_) );
	OAI21X1 OAI21X1_450 ( .A(_1743_), .B(_1754_), .C(_1752_), .Y(_1545_) );
	MUX2X1 MUX2X1_19 ( .A(ALU_op_1_), .B(_1747_), .S(ALU_op_0_), .Y(_1546_) );
	NAND2X1 NAND2X1_224 ( .A(ALU_BI_0_), .B(_1745_), .Y(_1547_) );
	NAND2X1 NAND2X1_225 ( .A(_1547_), .B(_1546_), .Y(_1548_) );
	AOI21X1 AOI21X1_129 ( .A(_1744_), .B(_1748_), .C(ALU_right), .Y(_1549_) );
	NAND2X1 NAND2X1_226 ( .A(_1549_), .B(_1548_), .Y(_1550_) );
	NAND3X1 NAND3X1_161 ( .A(_1751_), .B(_1753_), .C(_1550_), .Y(_1551_) );
	AOI21X1 AOI21X1_130 ( .A(_1545_), .B(_1551_), .C(_1742_), .Y(_1552_) );
	INVX1 INVX1_155 ( .A(_1742_), .Y(_1553_) );
	OAI21X1 OAI21X1_451 ( .A(_1752_), .B(_1754_), .C(_1545_), .Y(_1554_) );
	OAI21X1 OAI21X1_452 ( .A(_1553_), .B(_1554_), .C(RDY_bF_buf8), .Y(_1555_) );
	OAI21X1 OAI21X1_453 ( .A(_1552_), .B(_1555_), .C(_1740_), .Y(_1544__0_) );
	NAND2X1 NAND2X1_227 ( .A(ADD_1_), .B(_1717__bF_buf2), .Y(_1556_) );
	NOR2X1 NOR2X1_260 ( .A(_1754_), .B(_1752_), .Y(_1557_) );
	OAI21X1 OAI21X1_454 ( .A(_1553_), .B(_1557_), .C(_1545_), .Y(_1558_) );
	NOR2X1 NOR2X1_261 ( .A(ALU_op_1_), .B(_1722_), .Y(_1559_) );
	AND2X2 AND2X2_44 ( .A(_1722_), .B(ALU_BI_1_), .Y(_1560_) );
	INVX1 INVX1_156 ( .A(AI_1_), .Y(_1561_) );
	OAI21X1 OAI21X1_455 ( .A(_1720_), .B(_1561_), .C(ALU_BI_1_), .Y(_1562_) );
	OAI21X1 OAI21X1_456 ( .A(_1559_), .B(_1560_), .C(_1562_), .Y(_1563_) );
	NAND2X1 NAND2X1_228 ( .A(ALU_BI_1_), .B(_1722_), .Y(_1564_) );
	AOI21X1 AOI21X1_131 ( .A(_1564_), .B(_1561_), .C(ALU_right), .Y(_1565_) );
	AOI22X1 AOI22X1_52 ( .A(ALU_right), .B(AI_2_), .C(_1565_), .D(_1563_), .Y(_1566_) );
	OAI21X1 OAI21X1_457 ( .A(ALU_op_3_), .B(ALU_BI_1_), .C(_1729_), .Y(_1567_) );
	OAI21X1 OAI21X1_458 ( .A(ALU_BI_1_), .B(_1731_), .C(_1567_), .Y(_1568_) );
	OAI21X1 OAI21X1_459 ( .A(_1736_), .B(ALU_op_2_), .C(_1568_), .Y(_1569_) );
	MUX2X1 MUX2X1_20 ( .A(_1569_), .B(_1568_), .S(_1566_), .Y(_1570_) );
	NAND2X1 NAND2X1_229 ( .A(_1570_), .B(_1558_), .Y(_1571_) );
	OAI21X1 OAI21X1_460 ( .A(_1736_), .B(ALU_op_2_), .C(_1753_), .Y(_1572_) );
	AOI22X1 AOI22X1_53 ( .A(_1752_), .B(_1572_), .C(_1742_), .D(_1551_), .Y(_1573_) );
	INVX1 INVX1_157 ( .A(AI_2_), .Y(_1574_) );
	NAND2X1 NAND2X1_230 ( .A(ALU_op_1_), .B(AI_1_), .Y(_1575_) );
	AOI22X1 AOI22X1_54 ( .A(ALU_BI_1_), .B(_1575_), .C(_1721_), .D(_1564_), .Y(_1576_) );
	INVX1 INVX1_158 ( .A(_1565_), .Y(_1577_) );
	OAI22X1 OAI22X1_59 ( .A(_1726_), .B(_1574_), .C(_1576_), .D(_1577_), .Y(_1578_) );
	AND2X2 AND2X2_45 ( .A(_1578_), .B(_1568_), .Y(_1579_) );
	INVX1 INVX1_159 ( .A(_1743_), .Y(_1580_) );
	AOI21X1 AOI21X1_132 ( .A(_1580_), .B(_1568_), .C(_1578_), .Y(_1581_) );
	OAI21X1 OAI21X1_461 ( .A(_1581_), .B(_1579_), .C(_1573_), .Y(_1582_) );
	NAND2X1 NAND2X1_231 ( .A(_1571_), .B(_1582_), .Y(_1583_) );
	OAI21X1 OAI21X1_462 ( .A(_1717__bF_buf1), .B(_1583_), .C(_1556_), .Y(_1544__1_) );
	NAND2X1 NAND2X1_232 ( .A(ADD_2_), .B(_1717__bF_buf0), .Y(_1584_) );
	NAND2X1 NAND2X1_233 ( .A(_1568_), .B(_1578_), .Y(_1585_) );
	OAI21X1 OAI21X1_463 ( .A(_1581_), .B(_1573_), .C(_1585_), .Y(_1586_) );
	INVX1 INVX1_160 ( .A(AI_3_), .Y(_1587_) );
	INVX1 INVX1_161 ( .A(ALU_BI_2_), .Y(_1588_) );
	NOR2X1 NOR2X1_262 ( .A(ALU_op_0_), .B(_1588_), .Y(_1589_) );
	OAI21X1 OAI21X1_464 ( .A(_1720_), .B(_1574_), .C(ALU_BI_2_), .Y(_1590_) );
	OAI21X1 OAI21X1_465 ( .A(_1559_), .B(_1589_), .C(_1590_), .Y(_1591_) );
	OAI21X1 OAI21X1_466 ( .A(ALU_op_0_), .B(_1588_), .C(_1574_), .Y(_1592_) );
	NAND3X1 NAND3X1_162 ( .A(_1726_), .B(_1592_), .C(_1591_), .Y(_1593_) );
	OAI21X1 OAI21X1_467 ( .A(_1726_), .B(_1587_), .C(_1593_), .Y(_1594_) );
	OAI21X1 OAI21X1_468 ( .A(ALU_op_3_), .B(ALU_BI_2_), .C(_1729_), .Y(_1595_) );
	OAI21X1 OAI21X1_469 ( .A(ALU_BI_2_), .B(_1731_), .C(_1595_), .Y(_1596_) );
	NAND2X1 NAND2X1_234 ( .A(_1596_), .B(_1594_), .Y(_1597_) );
	NAND2X1 NAND2X1_235 ( .A(ALU_right), .B(AI_3_), .Y(_1598_) );
	OAI21X1 OAI21X1_470 ( .A(_1736_), .B(ALU_op_2_), .C(_1596_), .Y(_1599_) );
	NAND3X1 NAND3X1_163 ( .A(_1598_), .B(_1593_), .C(_1599_), .Y(_1600_) );
	AND2X2 AND2X2_46 ( .A(_1597_), .B(_1600_), .Y(_1601_) );
	NAND2X1 NAND2X1_236 ( .A(_1601_), .B(_1586_), .Y(_1602_) );
	NAND2X1 NAND2X1_237 ( .A(_1600_), .B(_1597_), .Y(_1603_) );
	NAND3X1 NAND3X1_164 ( .A(_1585_), .B(_1603_), .C(_1571_), .Y(_1604_) );
	NAND2X1 NAND2X1_238 ( .A(_1602_), .B(_1604_), .Y(_1605_) );
	OAI21X1 OAI21X1_471 ( .A(_1717__bF_buf3), .B(_1605_), .C(_1584_), .Y(_1544__2_) );
	NAND2X1 NAND2X1_239 ( .A(ADD_3_), .B(_1717__bF_buf2), .Y(_1606_) );
	AOI22X1 AOI22X1_55 ( .A(_1594_), .B(_1596_), .C(_1601_), .D(_1586_), .Y(_1607_) );
	INVX1 INVX1_162 ( .A(AI_4_), .Y(_1608_) );
	INVX1 INVX1_163 ( .A(ALU_BI_3_), .Y(_1609_) );
	NOR2X1 NOR2X1_263 ( .A(ALU_op_0_), .B(_1609_), .Y(_1610_) );
	OAI21X1 OAI21X1_472 ( .A(_1720_), .B(_1587_), .C(ALU_BI_3_), .Y(_1611_) );
	OAI21X1 OAI21X1_473 ( .A(_1559_), .B(_1610_), .C(_1611_), .Y(_1612_) );
	OAI21X1 OAI21X1_474 ( .A(ALU_op_0_), .B(_1609_), .C(_1587_), .Y(_1613_) );
	NAND3X1 NAND3X1_165 ( .A(_1726_), .B(_1613_), .C(_1612_), .Y(_1614_) );
	OAI21X1 OAI21X1_475 ( .A(_1726_), .B(_1608_), .C(_1614_), .Y(_1615_) );
	OAI21X1 OAI21X1_476 ( .A(ALU_op_3_), .B(ALU_BI_3_), .C(_1729_), .Y(_1616_) );
	OAI21X1 OAI21X1_477 ( .A(ALU_BI_3_), .B(_1731_), .C(_1616_), .Y(_1617_) );
	NAND2X1 NAND2X1_240 ( .A(_1617_), .B(_1615_), .Y(_1618_) );
	AND2X2 AND2X2_47 ( .A(_1617_), .B(_1580_), .Y(_1619_) );
	OAI21X1 OAI21X1_478 ( .A(_1615_), .B(_1619_), .C(_1618_), .Y(_1620_) );
	XNOR2X1 XNOR2X1_9 ( .A(_1607_), .B(_1620_), .Y(_1621_) );
	OAI21X1 OAI21X1_479 ( .A(_1717__bF_buf1), .B(_1621_), .C(_1606_), .Y(_1544__3_) );
	NAND2X1 NAND2X1_241 ( .A(ADD_4_), .B(_1717__bF_buf0), .Y(_1622_) );
	NAND3X1 NAND3X1_166 ( .A(_1585_), .B(_1601_), .C(_1571_), .Y(_1623_) );
	NAND2X1 NAND2X1_242 ( .A(_1603_), .B(_1586_), .Y(_1624_) );
	NAND3X1 NAND3X1_167 ( .A(_1624_), .B(_1583_), .C(_1623_), .Y(_1625_) );
	NAND2X1 NAND2X1_243 ( .A(ALU_BCD), .B(_1625_), .Y(_1626_) );
	NAND2X1 NAND2X1_244 ( .A(_1618_), .B(_1607_), .Y(_1627_) );
	OAI21X1 OAI21X1_480 ( .A(_1615_), .B(_1619_), .C(_1627_), .Y(_1628_) );
	OAI21X1 OAI21X1_481 ( .A(_1626_), .B(_1621_), .C(_1628_), .Y(_1629_) );
	NAND2X1 NAND2X1_245 ( .A(ALU_right), .B(AI_5_), .Y(_1630_) );
	AND2X2 AND2X2_48 ( .A(_1722_), .B(ALU_BI_4_), .Y(_1631_) );
	NAND2X1 NAND2X1_246 ( .A(AI_4_), .B(_1631_), .Y(_1632_) );
	AOI22X1 AOI22X1_56 ( .A(_1720_), .B(ALU_BI_4_), .C(_1721_), .D(_1632_), .Y(_1633_) );
	OAI21X1 OAI21X1_482 ( .A(AI_4_), .B(_1631_), .C(_1726_), .Y(_1634_) );
	OAI21X1 OAI21X1_483 ( .A(_1634_), .B(_1633_), .C(_1630_), .Y(_1635_) );
	NAND2X1 NAND2X1_247 ( .A(ALU_BI_4_), .B(_1733_), .Y(_1636_) );
	OAI21X1 OAI21X1_484 ( .A(ALU_BI_4_), .B(_1731_), .C(_1636_), .Y(_1637_) );
	OAI21X1 OAI21X1_485 ( .A(_1743_), .B(_1637_), .C(_1635_), .Y(_1638_) );
	OAI21X1 OAI21X1_486 ( .A(_1635_), .B(_1637_), .C(_1638_), .Y(_1639_) );
	INVX1 INVX1_164 ( .A(_1639_), .Y(_1640_) );
	NOR2X1 NOR2X1_264 ( .A(_1640_), .B(_1629_), .Y(_1641_) );
	OR2X2 OR2X2_33 ( .A(_1615_), .B(_1619_), .Y(_1642_) );
	XOR2X1 XOR2X1_2 ( .A(_1607_), .B(_1620_), .Y(_1643_) );
	INVX1 INVX1_165 ( .A(ALU_BCD), .Y(_1644_) );
	AOI21X1 AOI21X1_133 ( .A(_1605_), .B(_1583_), .C(_1644_), .Y(_1645_) );
	AOI22X1 AOI22X1_57 ( .A(_1642_), .B(_1627_), .C(_1643_), .D(_1645_), .Y(_1646_) );
	OAI21X1 OAI21X1_487 ( .A(_1639_), .B(_1646_), .C(RDY_bF_buf7), .Y(_1647_) );
	OAI21X1 OAI21X1_488 ( .A(_1641_), .B(_1647_), .C(_1622_), .Y(_1544__4_) );
	NAND2X1 NAND2X1_248 ( .A(ADD_5_), .B(_1717__bF_buf3), .Y(_1648_) );
	OAI21X1 OAI21X1_489 ( .A(_1639_), .B(_1646_), .C(_1638_), .Y(_1649_) );
	NAND2X1 NAND2X1_249 ( .A(ALU_right), .B(AI_6_), .Y(_1650_) );
	AND2X2 AND2X2_49 ( .A(_1722_), .B(ALU_BI_5_), .Y(_1651_) );
	NAND2X1 NAND2X1_250 ( .A(AI_5_), .B(_1651_), .Y(_1652_) );
	AOI22X1 AOI22X1_58 ( .A(_1720_), .B(ALU_BI_5_), .C(_1721_), .D(_1652_), .Y(_1653_) );
	OAI21X1 OAI21X1_490 ( .A(AI_5_), .B(_1651_), .C(_1726_), .Y(_1654_) );
	OAI21X1 OAI21X1_491 ( .A(_1654_), .B(_1653_), .C(_1650_), .Y(_1655_) );
	OAI21X1 OAI21X1_492 ( .A(ALU_op_3_), .B(ALU_BI_5_), .C(_1729_), .Y(_1656_) );
	OAI21X1 OAI21X1_493 ( .A(ALU_BI_5_), .B(_1731_), .C(_1656_), .Y(_1657_) );
	NAND2X1 NAND2X1_251 ( .A(_1657_), .B(_1655_), .Y(_1658_) );
	OAI21X1 OAI21X1_494 ( .A(_1736_), .B(ALU_op_2_), .C(_1657_), .Y(_1659_) );
	INVX1 INVX1_166 ( .A(_1659_), .Y(_1660_) );
	OAI21X1 OAI21X1_495 ( .A(_1655_), .B(_1660_), .C(_1658_), .Y(_1661_) );
	INVX1 INVX1_167 ( .A(_1661_), .Y(_1662_) );
	NAND2X1 NAND2X1_252 ( .A(_1662_), .B(_1649_), .Y(_1663_) );
	INVX1 INVX1_168 ( .A(_1637_), .Y(_1664_) );
	OAI21X1 OAI21X1_496 ( .A(_1736_), .B(ALU_op_2_), .C(_1664_), .Y(_1665_) );
	AOI22X1 AOI22X1_59 ( .A(_1635_), .B(_1665_), .C(_1640_), .D(_1629_), .Y(_1666_) );
	NAND2X1 NAND2X1_253 ( .A(_1661_), .B(_1666_), .Y(_1667_) );
	NAND2X1 NAND2X1_254 ( .A(_1667_), .B(_1663_), .Y(_1668_) );
	OAI21X1 OAI21X1_497 ( .A(_1717__bF_buf2), .B(_1668_), .C(_1648_), .Y(_1544__5_) );
	NAND2X1 NAND2X1_255 ( .A(ADD_6_), .B(_1717__bF_buf1), .Y(_1669_) );
	OAI21X1 OAI21X1_498 ( .A(_1661_), .B(_1666_), .C(_1658_), .Y(_1670_) );
	AND2X2 AND2X2_50 ( .A(_1722_), .B(ALU_BI_6_), .Y(_1671_) );
	NAND2X1 NAND2X1_256 ( .A(AI_6_), .B(_1671_), .Y(_1672_) );
	AOI22X1 AOI22X1_60 ( .A(_1720_), .B(ALU_BI_6_), .C(_1721_), .D(_1672_), .Y(_1673_) );
	OAI21X1 OAI21X1_499 ( .A(AI_6_), .B(_1671_), .C(_1726_), .Y(_1674_) );
	OAI22X1 OAI22X1_60 ( .A(_1716_), .B(_1726_), .C(_1674_), .D(_1673_), .Y(_1675_) );
	INVX1 INVX1_169 ( .A(_1733_), .Y(_1676_) );
	OAI21X1 OAI21X1_500 ( .A(ALU_op_3_), .B(ALU_BI_6_), .C(ALU_op_2_), .Y(_1677_) );
	OAI21X1 OAI21X1_501 ( .A(ALU_BI_6_), .B(_1676_), .C(_1677_), .Y(_1678_) );
	INVX1 INVX1_170 ( .A(_1678_), .Y(_1679_) );
	NAND2X1 NAND2X1_257 ( .A(_1679_), .B(_1675_), .Y(_1680_) );
	NOR2X1 NOR2X1_265 ( .A(ALU_op_3_), .B(_1678_), .Y(_1681_) );
	OAI21X1 OAI21X1_502 ( .A(_1675_), .B(_1681_), .C(_1680_), .Y(_1682_) );
	INVX1 INVX1_171 ( .A(_1682_), .Y(_1683_) );
	NAND2X1 NAND2X1_258 ( .A(_1683_), .B(_1670_), .Y(_1684_) );
	NAND3X1 NAND3X1_168 ( .A(_1658_), .B(_1682_), .C(_1663_), .Y(_1685_) );
	NAND2X1 NAND2X1_259 ( .A(_1685_), .B(_1684_), .Y(_1686_) );
	OAI21X1 OAI21X1_503 ( .A(_1717__bF_buf0), .B(_1686_), .C(_1669_), .Y(_1544__6_) );
	INVX1 INVX1_172 ( .A(ADD_7_), .Y(_1687_) );
	AOI22X1 AOI22X1_61 ( .A(_1655_), .B(_1657_), .C(_1662_), .D(_1649_), .Y(_1688_) );
	OAI21X1 OAI21X1_504 ( .A(_1682_), .B(_1688_), .C(_1680_), .Y(_1689_) );
	OAI21X1 OAI21X1_505 ( .A(_1743_), .B(_1735_), .C(_1728_), .Y(_1690_) );
	OAI21X1 OAI21X1_506 ( .A(_1728_), .B(_1735_), .C(_1690_), .Y(_1691_) );
	NAND2X1 NAND2X1_260 ( .A(_1691_), .B(_1689_), .Y(_1692_) );
	INVX1 INVX1_173 ( .A(_1691_), .Y(_1693_) );
	NAND3X1 NAND3X1_169 ( .A(_1680_), .B(_1693_), .C(_1684_), .Y(_1694_) );
	NAND2X1 NAND2X1_261 ( .A(_1694_), .B(_1692_), .Y(_1695_) );
	NAND2X1 NAND2X1_262 ( .A(RDY_bF_buf6), .B(_1695_), .Y(_1696_) );
	OAI21X1 OAI21X1_507 ( .A(_1687_), .B(RDY_bF_buf5), .C(_1696_), .Y(_1544__7_) );
	NAND2X1 NAND2X1_263 ( .A(ALU_HC), .B(_1717__bF_buf3), .Y(_1697_) );
	OAI21X1 OAI21X1_508 ( .A(_1717__bF_buf2), .B(_1646_), .C(_1697_), .Y(_1542_) );
	INVX1 INVX1_174 ( .A(ALU_N), .Y(_1698_) );
	OAI21X1 OAI21X1_509 ( .A(RDY_bF_buf4), .B(_1698_), .C(_1696_), .Y(_1543_) );
	NOR2X1 NOR2X1_266 ( .A(_1726_), .B(_1748_), .Y(_1699_) );
	INVX1 INVX1_175 ( .A(_1680_), .Y(_1700_) );
	AOI22X1 AOI22X1_62 ( .A(_1728_), .B(_1737_), .C(_1700_), .D(_1693_), .Y(_1701_) );
	NAND2X1 NAND2X1_264 ( .A(_1683_), .B(_1693_), .Y(_1702_) );
	OAI21X1 OAI21X1_510 ( .A(_1702_), .B(_1688_), .C(_1701_), .Y(_1703_) );
	NAND2X1 NAND2X1_265 ( .A(_1699_), .B(_1703_), .Y(_1704_) );
	OR2X2 OR2X2_34 ( .A(_1703_), .B(_1699_), .Y(_1705_) );
	AOI21X1 AOI21X1_134 ( .A(_1686_), .B(_1668_), .C(_1644_), .Y(_1706_) );
	AOI22X1 AOI22X1_63 ( .A(_1704_), .B(_1705_), .C(_1695_), .D(_1706_), .Y(_1707_) );
	NAND2X1 NAND2X1_266 ( .A(ALU_CO), .B(_1717__bF_buf1), .Y(_1708_) );
	OAI21X1 OAI21X1_511 ( .A(_1717__bF_buf0), .B(_1707_), .C(_1708_), .Y(_1541_) );
	XOR2X1 XOR2X1_3 ( .A(ALU_AI7), .B(ALU_BI7), .Y(_1709_) );
	XNOR2X1 XNOR2X1_10 ( .A(ALU_N), .B(ALU_CO), .Y(_1710_) );
	XNOR2X1 XNOR2X1_11 ( .A(_1709_), .B(_1710_), .Y(ALU_V) );
	DFFPOSX1 DFFPOSX1_126 ( .CLK(clk_bF_buf0), .D(_1541_), .Q(ALU_CO) );
	DFFPOSX1 DFFPOSX1_127 ( .CLK(clk_bF_buf11), .D(_1543_), .Q(ALU_N) );
	DFFPOSX1 DFFPOSX1_128 ( .CLK(clk_bF_buf10), .D(_1542_), .Q(ALU_HC) );
	DFFPOSX1 DFFPOSX1_129 ( .CLK(clk_bF_buf9), .D(_1544__0_), .Q(ADD_0_) );
	DFFPOSX1 DFFPOSX1_130 ( .CLK(clk_bF_buf8), .D(_1544__1_), .Q(ADD_1_) );
	DFFPOSX1 DFFPOSX1_131 ( .CLK(clk_bF_buf7), .D(_1544__2_), .Q(ADD_2_) );
	DFFPOSX1 DFFPOSX1_132 ( .CLK(clk_bF_buf6), .D(_1544__3_), .Q(ADD_3_) );
	DFFPOSX1 DFFPOSX1_133 ( .CLK(clk_bF_buf5), .D(_1544__4_), .Q(ADD_4_) );
	DFFPOSX1 DFFPOSX1_134 ( .CLK(clk_bF_buf4), .D(_1544__5_), .Q(ADD_5_) );
	DFFPOSX1 DFFPOSX1_135 ( .CLK(clk_bF_buf3), .D(_1544__6_), .Q(ADD_6_) );
	DFFPOSX1 DFFPOSX1_136 ( .CLK(clk_bF_buf2), .D(_1544__7_), .Q(ADD_7_) );
	DFFPOSX1 DFFPOSX1_137 ( .CLK(clk_bF_buf1), .D(_1540_), .Q(ALU_BI7) );
	DFFPOSX1 DFFPOSX1_138 ( .CLK(clk_bF_buf0), .D(_1539_), .Q(ALU_AI7) );
endmodule
