module pic27ch ( gnd, vdd, in4, in17, in30, in43, in56, in69, in82, in95, in108, in1, in11, in24, in37, in50, in63, in76, in89, in102, in8, in21, in34, in47, in60, in73, in86, in99, in112, in14, in27, in40, in53, in66, in79, in92, in105, in115, out223, out329, out370, out421, out430, out431, out432);

input gnd, vdd;
input in4;
input in17;
input in30;
input in43;
input in56;
input in69;
input in82;
input in95;
input in108;
input in1;
input in11;
input in24;
input in37;
input in50;
input in63;
input in76;
input in89;
input in102;
input in8;
input in21;
input in34;
input in47;
input in60;
input in73;
input in86;
input in99;
input in112;
input in14;
input in27;
input in40;
input in53;
input in66;
input in79;
input in92;
input in105;
input in115;
output out223;
output out329;
output out370;
output out421;
output out430;
output out431;
output out432;

BUFX4 BUFX4_1 ( .gnd(gnd), .vdd(vdd), .A(_1_), .Y(_1__bF_buf3) );
BUFX4 BUFX4_2 ( .gnd(gnd), .vdd(vdd), .A(_1_), .Y(_1__bF_buf2) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_1_), .Y(_1__bF_buf1) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_1_), .Y(_1__bF_buf0) );
BUFX4 BUFX4_3 ( .gnd(gnd), .vdd(vdd), .A(_0_), .Y(_0__bF_buf3) );
BUFX4 BUFX4_4 ( .gnd(gnd), .vdd(vdd), .A(_0_), .Y(_0__bF_buf2) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_0_), .Y(_0__bF_buf1) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_0_), .Y(_0__bF_buf0) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_0__bF_buf0), .Y(out223) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_1__bF_buf3), .Y(out329) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_2_), .Y(out370) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_3_), .Y(out421) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_4_), .Y(out430) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_5_), .Y(out431) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_6_), .Y(out432) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(in102), .Y(_7_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(in108), .B(_7_), .Y(_8_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(in82), .Y(_9_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(in95), .Y(_10_) );
OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(in76), .B(_9_), .C(_10_), .D(in89), .Y(_11_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(in56), .Y(_12_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(in69), .Y(_13_) );
OAI22X1 OAI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(in50), .B(_12_), .C(_13_), .D(in63), .Y(_14_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_11_), .B(_14_), .Y(_15_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(in30), .Y(_16_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(in43), .Y(_17_) );
OAI22X1 OAI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(in24), .B(_16_), .C(_17_), .D(in37), .Y(_18_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(in4), .Y(_19_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(in17), .Y(_20_) );
OAI22X1 OAI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(in1), .B(_19_), .C(_20_), .D(in11), .Y(_21_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_18_), .B(_21_), .Y(_22_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(_15_), .C(_22_), .Y(_0_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_15_), .B(_22_), .Y(_23_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(_23_), .Y(Ckt432_M1_X1_0_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_10_), .B(in89), .Y(_24_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_24_), .B(_0__bF_buf3), .Y(Ckt432_M1_X1_1_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_9_), .B(in76), .Y(_25_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_25_), .B(_0__bF_buf3), .Y(Ckt432_M1_X1_2_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_13_), .B(in63), .Y(_26_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_0__bF_buf3), .Y(Ckt432_M1_X1_3_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(in50), .Y(_27_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_27_), .B(_0__bF_buf2), .Y(Ckt432_M1_X1_4_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_17_), .B(in37), .Y(_28_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_28_), .B(_0__bF_buf1), .Y(Ckt432_M1_X1_5_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_16_), .B(in24), .Y(_29_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_29_), .B(_0__bF_buf1), .Y(Ckt432_M1_X1_6_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(in11), .Y(_30_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_30_), .B(_0__bF_buf0), .Y(Ckt432_M1_X1_7_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(_19_), .B(in1), .Y(_31_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_31_), .B(_0__bF_buf2), .Y(Ckt432_M1_X1_8_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(in112), .Y(_32_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(in108), .B(Ckt432_M1_X1_0_), .C(_32_), .Y(_33_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(in4), .B(Ckt432_M1_X1_8_), .Y(_34_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(in17), .B(Ckt432_M1_X1_7_), .Y(_35_) );
OAI22X1 OAI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(in8), .B(_34_), .C(in21), .D(_35_), .Y(_36_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(Ckt432_M1_X1_6_), .B(in30), .Y(_37_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(Ckt432_M1_X1_5_), .B(in43), .Y(_38_) );
OAI22X1 OAI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(in34), .B(_37_), .C(in47), .D(_38_), .Y(_39_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_36_), .B(_39_), .Y(_40_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(Ckt432_M1_X1_2_), .B(in82), .Y(_41_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(Ckt432_M1_X1_1_), .B(in95), .Y(_42_) );
OAI22X1 OAI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(in86), .B(_41_), .C(in99), .D(_42_), .Y(_43_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(Ckt432_M1_X1_4_), .B(in56), .Y(_44_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(Ckt432_M1_X1_3_), .B(in69), .Y(_45_) );
OAI22X1 OAI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(in60), .B(_44_), .C(in73), .D(_45_), .Y(_46_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_43_), .B(_46_), .Y(_47_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_33_), .B(_40_), .C(_47_), .Y(_1_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_47_), .Y(_48_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_33_), .B(_48_), .Y(Ckt432_M2_X2_0_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_42_), .B(in99), .Y(_49_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_49_), .B(_1__bF_buf3), .Y(Ckt432_M2_X2_1_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_41_), .B(in86), .Y(_50_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_50_), .B(_1__bF_buf3), .Y(Ckt432_M2_X2_2_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_45_), .B(in73), .Y(_51_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_51_), .B(_1__bF_buf0), .Y(Ckt432_M2_X2_3_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_44_), .B(in60), .Y(_52_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(_1__bF_buf0), .Y(Ckt432_M2_X2_4_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(_38_), .B(in47), .Y(_53_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_53_), .B(_1__bF_buf1), .Y(Ckt432_M2_X2_5_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(_37_), .B(in34), .Y(_54_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_54_), .B(_1__bF_buf1), .Y(Ckt432_M2_X2_6_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(_35_), .B(in21), .Y(_55_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_55_), .B(_1__bF_buf2), .Y(Ckt432_M2_X2_7_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(_34_), .B(in8), .Y(_56_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_56_), .B(_1__bF_buf2), .Y(Ckt432_M2_X2_8_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(Ckt432_M2_X2_5_), .B(Ckt432_M1_X1_5_), .Y(_57_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(in53), .Y(_58_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(in43), .B(_58_), .Y(_59_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(Ckt432_M1_X1_6_), .B(in30), .Y(_60_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(in40), .Y(_61_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(Ckt432_M2_X2_6_), .B(_61_), .Y(_62_) );
OAI22X1 OAI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(_57_), .B(_59_), .C(_60_), .D(_62_), .Y(_63_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(Ckt432_M1_X1_1_), .B(in95), .Y(_64_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(Ckt432_M2_X2_1_), .Y(_65_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(in105), .B(_65_), .Y(_66_) );
AOI21X1 AOI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_64_), .B(_66_), .C(_63_), .Y(_67_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(Ckt432_M2_X2_7_), .B(Ckt432_M1_X1_7_), .Y(_68_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(in17), .Y(_69_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(in27), .B(_69_), .Y(_70_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(Ckt432_M2_X2_4_), .B(Ckt432_M1_X1_4_), .Y(_71_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(in56), .Y(_72_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(in66), .B(_72_), .Y(_73_) );
AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_70_), .B(_68_), .C(_71_), .D(_73_), .Y(_74_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(Ckt432_M2_X2_0_), .B(Ckt432_M1_X1_0_), .Y(_75_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(in115), .Y(_76_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(in108), .B(_76_), .Y(_77_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(Ckt432_M1_X1_3_), .B(in69), .Y(_78_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(in79), .Y(_79_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(Ckt432_M2_X2_3_), .B(_79_), .Y(_80_) );
OAI22X1 OAI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_75_), .B(_77_), .C(_78_), .D(_80_), .Y(_81_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(Ckt432_M2_X2_8_), .B(Ckt432_M1_X1_8_), .Y(_82_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(in14), .Y(_83_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(in4), .B(_83_), .Y(_84_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(Ckt432_M1_X1_2_), .B(in82), .Y(_85_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(in92), .Y(_86_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(Ckt432_M2_X2_2_), .B(_86_), .Y(_87_) );
OAI22X1 OAI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(_82_), .B(_84_), .C(_85_), .D(_87_), .Y(_88_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_81_), .B(_88_), .Y(_89_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_74_), .B(_67_), .C(_89_), .Y(_2_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_2_), .B(in115), .Y(_90_) );
AOI22X1 AOI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_0__bF_buf2), .B(in102), .C(_1__bF_buf2), .D(in112), .Y(_91_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(in108), .B(_90_), .C(_91_), .Y(Ckt432_I_0_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_2_), .B(in105), .Y(_92_) );
AOI22X1 AOI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_0__bF_buf3), .B(in89), .C(_1__bF_buf3), .D(in99), .Y(_93_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(in95), .B(_92_), .C(_93_), .Y(Ckt432_I_1_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_2_), .B(in92), .Y(_94_) );
AOI22X1 AOI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_0__bF_buf3), .B(in76), .C(_1__bF_buf3), .D(in86), .Y(_95_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(in82), .B(_94_), .C(_95_), .Y(Ckt432_I_2_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_2_), .B(in79), .Y(_96_) );
AOI22X1 AOI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_0__bF_buf2), .B(in63), .C(_1__bF_buf0), .D(in73), .Y(_97_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(in69), .B(_96_), .C(_97_), .Y(Ckt432_I_3_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_2_), .B(in66), .Y(_98_) );
AOI22X1 AOI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_0__bF_buf2), .B(in50), .C(_1__bF_buf0), .D(in60), .Y(_99_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(in56), .B(_98_), .C(_99_), .Y(Ckt432_I_4_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_2_), .B(in53), .Y(_100_) );
AOI22X1 AOI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_0__bF_buf1), .B(in37), .C(_1__bF_buf1), .D(in47), .Y(_101_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(in43), .B(_100_), .C(_101_), .Y(Ckt432_I_5_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_2_), .B(in40), .Y(_102_) );
AOI22X1 AOI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_0__bF_buf1), .B(in24), .C(_1__bF_buf1), .D(in34), .Y(_103_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(in30), .B(_102_), .C(_103_), .Y(Ckt432_I_6_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_2_), .B(in27), .Y(_104_) );
AOI22X1 AOI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(_0__bF_buf0), .B(in11), .C(_1__bF_buf2), .D(in21), .Y(_105_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(in17), .B(_104_), .C(_105_), .Y(Ckt432_I_7_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_2_), .B(in14), .Y(_106_) );
AOI22X1 AOI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_0__bF_buf0), .B(in1), .C(_1__bF_buf2), .D(in8), .Y(_107_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(in4), .B(_106_), .C(_107_), .Y(Ckt432_I_8_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(Ckt432_I_8_), .Y(_108_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(Ckt432_I_4_), .B(Ckt432_I_5_), .Y(_109_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(Ckt432_I_6_), .B(Ckt432_I_7_), .Y(_110_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_109_), .B(_110_), .Y(_111_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(Ckt432_I_2_), .B(Ckt432_I_3_), .Y(_112_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(Ckt432_I_0_), .B(Ckt432_I_1_), .Y(_113_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_112_), .B(_113_), .Y(_114_) );
AOI21X1 AOI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_111_), .B(_114_), .C(_108_), .Y(_3_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(_111_), .Y(_4_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(Ckt432_I_3_), .Y(_115_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(Ckt432_I_6_), .B(_115_), .C(_109_), .Y(_116_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(Ckt432_I_2_), .Y(_117_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_117_), .B(_109_), .Y(_118_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_110_), .B(_118_), .C(_116_), .Y(_5_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(Ckt432_I_1_), .B(_117_), .C(Ckt432_I_5_), .Y(_119_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(Ckt432_I_6_), .B(_119_), .Y(_120_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(Ckt432_I_7_), .B(_116_), .C(_120_), .Y(_6_) );
endmodule
